// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Feb 19 2025 16:49:25

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "LED_Blink_Top_Module" view "INTERFACE"

module LED_Blink_Top_Module (
    o_LED_3,
    o_LED_1,
    i_Clk,
    o_LED_4,
    o_LED_2);

    output o_LED_3;
    output o_LED_1;
    input i_Clk;
    output o_LED_4;
    output o_LED_2;

    wire N__4823;
    wire N__4822;
    wire N__4821;
    wire N__4812;
    wire N__4811;
    wire N__4810;
    wire N__4803;
    wire N__4802;
    wire N__4801;
    wire N__4794;
    wire N__4793;
    wire N__4792;
    wire N__4785;
    wire N__4784;
    wire N__4783;
    wire N__4766;
    wire N__4763;
    wire N__4760;
    wire N__4757;
    wire N__4756;
    wire N__4753;
    wire N__4750;
    wire N__4747;
    wire N__4742;
    wire N__4741;
    wire N__4738;
    wire N__4735;
    wire N__4730;
    wire N__4729;
    wire N__4726;
    wire N__4723;
    wire N__4718;
    wire N__4715;
    wire N__4714;
    wire N__4709;
    wire N__4706;
    wire N__4703;
    wire N__4702;
    wire N__4699;
    wire N__4696;
    wire N__4691;
    wire N__4688;
    wire N__4685;
    wire N__4682;
    wire N__4679;
    wire N__4678;
    wire N__4675;
    wire N__4672;
    wire N__4667;
    wire N__4664;
    wire N__4661;
    wire N__4660;
    wire N__4657;
    wire N__4654;
    wire N__4649;
    wire N__4648;
    wire N__4647;
    wire N__4646;
    wire N__4645;
    wire N__4644;
    wire N__4643;
    wire N__4642;
    wire N__4641;
    wire N__4640;
    wire N__4639;
    wire N__4638;
    wire N__4637;
    wire N__4636;
    wire N__4629;
    wire N__4626;
    wire N__4617;
    wire N__4614;
    wire N__4603;
    wire N__4592;
    wire N__4591;
    wire N__4590;
    wire N__4587;
    wire N__4586;
    wire N__4585;
    wire N__4584;
    wire N__4581;
    wire N__4580;
    wire N__4579;
    wire N__4578;
    wire N__4575;
    wire N__4574;
    wire N__4573;
    wire N__4572;
    wire N__4571;
    wire N__4570;
    wire N__4563;
    wire N__4552;
    wire N__4541;
    wire N__4538;
    wire N__4529;
    wire N__4528;
    wire N__4525;
    wire N__4524;
    wire N__4521;
    wire N__4520;
    wire N__4519;
    wire N__4518;
    wire N__4517;
    wire N__4516;
    wire N__4515;
    wire N__4514;
    wire N__4513;
    wire N__4512;
    wire N__4511;
    wire N__4506;
    wire N__4499;
    wire N__4496;
    wire N__4489;
    wire N__4480;
    wire N__4475;
    wire N__4466;
    wire N__4463;
    wire N__4462;
    wire N__4459;
    wire N__4456;
    wire N__4453;
    wire N__4450;
    wire N__4445;
    wire N__4444;
    wire N__4443;
    wire N__4442;
    wire N__4441;
    wire N__4440;
    wire N__4439;
    wire N__4438;
    wire N__4437;
    wire N__4436;
    wire N__4435;
    wire N__4434;
    wire N__4433;
    wire N__4432;
    wire N__4431;
    wire N__4430;
    wire N__4429;
    wire N__4428;
    wire N__4427;
    wire N__4426;
    wire N__4425;
    wire N__4424;
    wire N__4423;
    wire N__4422;
    wire N__4373;
    wire N__4370;
    wire N__4367;
    wire N__4366;
    wire N__4363;
    wire N__4360;
    wire N__4355;
    wire N__4352;
    wire N__4349;
    wire N__4346;
    wire N__4343;
    wire N__4340;
    wire N__4337;
    wire N__4334;
    wire N__4333;
    wire N__4330;
    wire N__4327;
    wire N__4322;
    wire N__4319;
    wire N__4316;
    wire N__4313;
    wire N__4310;
    wire N__4309;
    wire N__4306;
    wire N__4303;
    wire N__4298;
    wire N__4295;
    wire N__4292;
    wire N__4289;
    wire N__4286;
    wire N__4283;
    wire N__4280;
    wire N__4277;
    wire N__4276;
    wire N__4273;
    wire N__4270;
    wire N__4265;
    wire N__4262;
    wire N__4259;
    wire N__4256;
    wire N__4253;
    wire N__4252;
    wire N__4249;
    wire N__4246;
    wire N__4241;
    wire N__4238;
    wire N__4235;
    wire N__4232;
    wire N__4231;
    wire N__4228;
    wire N__4225;
    wire N__4220;
    wire N__4217;
    wire N__4214;
    wire N__4211;
    wire N__4208;
    wire N__4205;
    wire N__4204;
    wire N__4201;
    wire N__4198;
    wire N__4193;
    wire N__4190;
    wire N__4189;
    wire N__4186;
    wire N__4183;
    wire N__4178;
    wire N__4175;
    wire N__4174;
    wire N__4171;
    wire N__4168;
    wire N__4163;
    wire N__4160;
    wire N__4157;
    wire N__4156;
    wire N__4153;
    wire N__4150;
    wire N__4145;
    wire N__4142;
    wire N__4139;
    wire N__4136;
    wire N__4135;
    wire N__4132;
    wire N__4129;
    wire N__4124;
    wire N__4121;
    wire N__4118;
    wire N__4115;
    wire N__4112;
    wire N__4109;
    wire N__4108;
    wire N__4105;
    wire N__4102;
    wire N__4097;
    wire N__4094;
    wire N__4091;
    wire N__4088;
    wire N__4085;
    wire N__4084;
    wire N__4081;
    wire N__4078;
    wire N__4073;
    wire N__4072;
    wire N__4069;
    wire N__4066;
    wire N__4063;
    wire N__4058;
    wire N__4057;
    wire N__4054;
    wire N__4051;
    wire N__4046;
    wire N__4045;
    wire N__4042;
    wire N__4039;
    wire N__4034;
    wire N__4033;
    wire N__4032;
    wire N__4029;
    wire N__4026;
    wire N__4023;
    wire N__4016;
    wire N__4013;
    wire N__4010;
    wire N__4007;
    wire N__4006;
    wire N__4003;
    wire N__4000;
    wire N__3995;
    wire N__3994;
    wire N__3991;
    wire N__3988;
    wire N__3983;
    wire N__3980;
    wire N__3977;
    wire N__3974;
    wire N__3971;
    wire N__3968;
    wire N__3965;
    wire N__3962;
    wire N__3961;
    wire N__3958;
    wire N__3955;
    wire N__3950;
    wire N__3949;
    wire N__3948;
    wire N__3947;
    wire N__3946;
    wire N__3945;
    wire N__3942;
    wire N__3941;
    wire N__3940;
    wire N__3939;
    wire N__3936;
    wire N__3933;
    wire N__3932;
    wire N__3929;
    wire N__3926;
    wire N__3921;
    wire N__3918;
    wire N__3909;
    wire N__3902;
    wire N__3893;
    wire N__3892;
    wire N__3889;
    wire N__3886;
    wire N__3885;
    wire N__3884;
    wire N__3883;
    wire N__3882;
    wire N__3881;
    wire N__3880;
    wire N__3879;
    wire N__3878;
    wire N__3871;
    wire N__3868;
    wire N__3865;
    wire N__3862;
    wire N__3857;
    wire N__3852;
    wire N__3847;
    wire N__3836;
    wire N__3835;
    wire N__3834;
    wire N__3833;
    wire N__3832;
    wire N__3831;
    wire N__3830;
    wire N__3829;
    wire N__3828;
    wire N__3825;
    wire N__3820;
    wire N__3815;
    wire N__3806;
    wire N__3797;
    wire N__3796;
    wire N__3793;
    wire N__3790;
    wire N__3787;
    wire N__3782;
    wire N__3781;
    wire N__3780;
    wire N__3777;
    wire N__3774;
    wire N__3771;
    wire N__3764;
    wire N__3763;
    wire N__3762;
    wire N__3761;
    wire N__3758;
    wire N__3755;
    wire N__3750;
    wire N__3747;
    wire N__3740;
    wire N__3739;
    wire N__3736;
    wire N__3733;
    wire N__3728;
    wire N__3725;
    wire N__3724;
    wire N__3721;
    wire N__3718;
    wire N__3713;
    wire N__3710;
    wire N__3707;
    wire N__3704;
    wire N__3703;
    wire N__3700;
    wire N__3697;
    wire N__3692;
    wire N__3691;
    wire N__3688;
    wire N__3685;
    wire N__3680;
    wire N__3679;
    wire N__3678;
    wire N__3677;
    wire N__3674;
    wire N__3667;
    wire N__3664;
    wire N__3659;
    wire N__3658;
    wire N__3655;
    wire N__3652;
    wire N__3647;
    wire N__3644;
    wire N__3641;
    wire N__3640;
    wire N__3637;
    wire N__3634;
    wire N__3629;
    wire N__3626;
    wire N__3623;
    wire N__3620;
    wire N__3617;
    wire N__3616;
    wire N__3613;
    wire N__3610;
    wire N__3605;
    wire N__3604;
    wire N__3601;
    wire N__3598;
    wire N__3593;
    wire N__3590;
    wire N__3589;
    wire N__3586;
    wire N__3583;
    wire N__3578;
    wire N__3577;
    wire N__3574;
    wire N__3571;
    wire N__3566;
    wire N__3563;
    wire N__3560;
    wire N__3557;
    wire N__3554;
    wire N__3551;
    wire N__3548;
    wire N__3545;
    wire N__3542;
    wire N__3539;
    wire N__3536;
    wire N__3533;
    wire N__3530;
    wire N__3529;
    wire N__3524;
    wire N__3521;
    wire N__3518;
    wire N__3515;
    wire N__3512;
    wire N__3509;
    wire N__3506;
    wire N__3503;
    wire N__3500;
    wire N__3497;
    wire N__3496;
    wire N__3491;
    wire N__3488;
    wire N__3485;
    wire N__3484;
    wire N__3479;
    wire N__3476;
    wire N__3475;
    wire N__3470;
    wire N__3467;
    wire N__3464;
    wire N__3461;
    wire N__3458;
    wire N__3455;
    wire N__3452;
    wire N__3449;
    wire N__3446;
    wire N__3443;
    wire N__3440;
    wire N__3437;
    wire N__3434;
    wire N__3431;
    wire N__3428;
    wire N__3427;
    wire N__3426;
    wire N__3425;
    wire N__3424;
    wire N__3423;
    wire N__3422;
    wire N__3421;
    wire N__3420;
    wire N__3419;
    wire N__3418;
    wire N__3415;
    wire N__3406;
    wire N__3397;
    wire N__3392;
    wire N__3383;
    wire N__3380;
    wire N__3377;
    wire N__3376;
    wire N__3375;
    wire N__3374;
    wire N__3373;
    wire N__3372;
    wire N__3371;
    wire N__3370;
    wire N__3369;
    wire N__3366;
    wire N__3363;
    wire N__3360;
    wire N__3357;
    wire N__3354;
    wire N__3351;
    wire N__3350;
    wire N__3347;
    wire N__3346;
    wire N__3345;
    wire N__3342;
    wire N__3339;
    wire N__3334;
    wire N__3329;
    wire N__3326;
    wire N__3321;
    wire N__3318;
    wire N__3311;
    wire N__3308;
    wire N__3303;
    wire N__3296;
    wire N__3287;
    wire N__3286;
    wire N__3285;
    wire N__3284;
    wire N__3283;
    wire N__3282;
    wire N__3281;
    wire N__3280;
    wire N__3279;
    wire N__3270;
    wire N__3269;
    wire N__3268;
    wire N__3265;
    wire N__3256;
    wire N__3253;
    wire N__3248;
    wire N__3239;
    wire N__3238;
    wire N__3235;
    wire N__3232;
    wire N__3227;
    wire N__3226;
    wire N__3223;
    wire N__3220;
    wire N__3215;
    wire N__3214;
    wire N__3211;
    wire N__3208;
    wire N__3205;
    wire N__3200;
    wire N__3199;
    wire N__3196;
    wire N__3193;
    wire N__3188;
    wire N__3185;
    wire N__3182;
    wire N__3179;
    wire N__3176;
    wire N__3173;
    wire N__3172;
    wire N__3171;
    wire N__3166;
    wire N__3163;
    wire N__3158;
    wire N__3155;
    wire N__3152;
    wire N__3149;
    wire N__3148;
    wire N__3145;
    wire N__3142;
    wire N__3137;
    wire N__3134;
    wire N__3131;
    wire N__3128;
    wire N__3125;
    wire N__3122;
    wire N__3119;
    wire N__3116;
    wire N__3113;
    wire N__3110;
    wire N__3109;
    wire N__3106;
    wire N__3103;
    wire N__3098;
    wire N__3097;
    wire N__3094;
    wire N__3091;
    wire N__3086;
    wire N__3085;
    wire N__3082;
    wire N__3079;
    wire N__3074;
    wire N__3071;
    wire N__3070;
    wire N__3067;
    wire N__3064;
    wire N__3061;
    wire N__3056;
    wire N__3055;
    wire N__3052;
    wire N__3049;
    wire N__3044;
    wire N__3041;
    wire N__3038;
    wire N__3035;
    wire N__3032;
    wire N__3031;
    wire N__3028;
    wire N__3025;
    wire N__3020;
    wire N__3017;
    wire N__3014;
    wire N__3013;
    wire N__3010;
    wire N__3007;
    wire N__3002;
    wire N__2999;
    wire N__2996;
    wire N__2993;
    wire N__2990;
    wire N__2987;
    wire N__2986;
    wire N__2983;
    wire N__2980;
    wire N__2975;
    wire N__2972;
    wire N__2971;
    wire N__2968;
    wire N__2965;
    wire N__2960;
    wire N__2957;
    wire N__2956;
    wire N__2953;
    wire N__2950;
    wire N__2947;
    wire N__2944;
    wire N__2939;
    wire N__2936;
    wire N__2933;
    wire N__2930;
    wire N__2929;
    wire N__2926;
    wire N__2923;
    wire N__2920;
    wire N__2917;
    wire N__2912;
    wire N__2911;
    wire N__2908;
    wire N__2905;
    wire N__2900;
    wire N__2899;
    wire N__2896;
    wire N__2893;
    wire N__2888;
    wire N__2885;
    wire N__2884;
    wire N__2881;
    wire N__2878;
    wire N__2873;
    wire N__2872;
    wire N__2869;
    wire N__2866;
    wire N__2861;
    wire N__2860;
    wire N__2857;
    wire N__2856;
    wire N__2855;
    wire N__2852;
    wire N__2847;
    wire N__2844;
    wire N__2841;
    wire N__2834;
    wire N__2833;
    wire N__2830;
    wire N__2827;
    wire N__2822;
    wire N__2821;
    wire N__2818;
    wire N__2815;
    wire N__2810;
    wire N__2807;
    wire N__2806;
    wire N__2803;
    wire N__2800;
    wire N__2795;
    wire N__2792;
    wire N__2789;
    wire N__2786;
    wire N__2783;
    wire N__2780;
    wire N__2777;
    wire N__2774;
    wire N__2771;
    wire N__2768;
    wire N__2765;
    wire N__2762;
    wire N__2759;
    wire N__2756;
    wire N__2753;
    wire N__2750;
    wire N__2747;
    wire N__2744;
    wire N__2741;
    wire N__2738;
    wire N__2735;
    wire N__2734;
    wire N__2731;
    wire N__2728;
    wire N__2723;
    wire N__2720;
    wire N__2719;
    wire N__2718;
    wire N__2717;
    wire N__2714;
    wire N__2711;
    wire N__2706;
    wire N__2703;
    wire N__2696;
    wire N__2693;
    wire N__2690;
    wire N__2687;
    wire N__2684;
    wire N__2683;
    wire N__2680;
    wire N__2677;
    wire N__2672;
    wire N__2671;
    wire N__2668;
    wire N__2665;
    wire N__2660;
    wire N__2659;
    wire N__2656;
    wire N__2653;
    wire N__2648;
    wire N__2645;
    wire N__2644;
    wire N__2641;
    wire N__2638;
    wire N__2633;
    wire N__2632;
    wire N__2629;
    wire N__2626;
    wire N__2621;
    wire N__2620;
    wire N__2619;
    wire N__2618;
    wire N__2617;
    wire N__2616;
    wire N__2613;
    wire N__2612;
    wire N__2609;
    wire N__2606;
    wire N__2597;
    wire N__2596;
    wire N__2595;
    wire N__2592;
    wire N__2589;
    wire N__2586;
    wire N__2583;
    wire N__2578;
    wire N__2575;
    wire N__2564;
    wire N__2563;
    wire N__2562;
    wire N__2561;
    wire N__2560;
    wire N__2557;
    wire N__2556;
    wire N__2555;
    wire N__2552;
    wire N__2549;
    wire N__2548;
    wire N__2545;
    wire N__2544;
    wire N__2539;
    wire N__2530;
    wire N__2523;
    wire N__2516;
    wire N__2515;
    wire N__2514;
    wire N__2513;
    wire N__2504;
    wire N__2503;
    wire N__2502;
    wire N__2501;
    wire N__2500;
    wire N__2499;
    wire N__2498;
    wire N__2495;
    wire N__2486;
    wire N__2481;
    wire N__2474;
    wire N__2471;
    wire N__2468;
    wire N__2465;
    wire N__2464;
    wire N__2461;
    wire N__2458;
    wire N__2453;
    wire N__2450;
    wire N__2447;
    wire N__2444;
    wire N__2443;
    wire N__2440;
    wire N__2437;
    wire N__2432;
    wire N__2431;
    wire N__2428;
    wire N__2425;
    wire N__2420;
    wire N__2417;
    wire N__2416;
    wire N__2413;
    wire N__2410;
    wire N__2405;
    wire N__2404;
    wire N__2401;
    wire N__2398;
    wire N__2393;
    wire N__2392;
    wire N__2391;
    wire N__2386;
    wire N__2383;
    wire N__2378;
    wire N__2375;
    wire N__2372;
    wire N__2371;
    wire N__2368;
    wire N__2365;
    wire N__2360;
    wire N__2357;
    wire N__2356;
    wire N__2353;
    wire N__2350;
    wire N__2347;
    wire N__2344;
    wire N__2339;
    wire N__2336;
    wire N__2333;
    wire N__2332;
    wire N__2329;
    wire N__2326;
    wire N__2321;
    wire N__2320;
    wire N__2317;
    wire N__2314;
    wire N__2309;
    wire N__2308;
    wire N__2305;
    wire N__2302;
    wire N__2297;
    wire N__2296;
    wire N__2293;
    wire N__2290;
    wire N__2285;
    wire N__2282;
    wire N__2279;
    wire N__2276;
    wire N__2273;
    wire N__2270;
    wire N__2267;
    wire N__2264;
    wire N__2261;
    wire N__2258;
    wire N__2255;
    wire N__2252;
    wire N__2251;
    wire N__2246;
    wire N__2243;
    wire N__2242;
    wire N__2237;
    wire N__2234;
    wire N__2233;
    wire N__2230;
    wire N__2225;
    wire N__2222;
    wire N__2221;
    wire N__2218;
    wire N__2215;
    wire N__2210;
    wire N__2207;
    wire N__2204;
    wire N__2201;
    wire N__2198;
    wire N__2195;
    wire N__2192;
    wire N__2189;
    wire N__2186;
    wire N__2183;
    wire N__2180;
    wire N__2177;
    wire N__2174;
    wire N__2171;
    wire N__2168;
    wire N__2165;
    wire N__2162;
    wire N__2159;
    wire N__2156;
    wire N__2153;
    wire VCCG0;
    wire GNDG0;
    wire bfn_7_5_0_;
    wire \LED_Blink_Inst.un4_r_count_5hz_cry_1 ;
    wire \LED_Blink_Inst.un4_r_count_5hz_cry_2 ;
    wire \LED_Blink_Inst.un4_r_count_5hz_cry_3 ;
    wire \LED_Blink_Inst.un4_r_count_5hz_cry_4 ;
    wire \LED_Blink_Inst.un4_r_count_5hz_cry_5 ;
    wire \LED_Blink_Inst.un4_r_count_5hz_cry_6 ;
    wire \LED_Blink_Inst.un4_r_count_5hz_cry_7 ;
    wire \LED_Blink_Inst.un4_r_count_5hz_cry_8 ;
    wire bfn_7_6_0_;
    wire \LED_Blink_Inst.un4_r_count_5hz_cry_9 ;
    wire \LED_Blink_Inst.un4_r_count_5hz_cry_10 ;
    wire \LED_Blink_Inst.un4_r_count_5hz_cry_11 ;
    wire \LED_Blink_Inst.un4_r_count_5hz_cry_12 ;
    wire \LED_Blink_Inst.un4_r_count_5hz_cry_13 ;
    wire \LED_Blink_Inst.un4_r_count_5hz_cry_14 ;
    wire \LED_Blink_Inst.un4_r_count_5hz_cry_15 ;
    wire \LED_Blink_Inst.un4_r_count_5hz_cry_16 ;
    wire bfn_7_7_0_;
    wire \LED_Blink_Inst.un4_r_count_5hz_cry_17 ;
    wire \LED_Blink_Inst.un4_r_count_5hz_cry_18 ;
    wire \LED_Blink_Inst.un4_r_count_5hz_cry_19 ;
    wire \LED_Blink_Inst.un4_r_count_5hz_cry_20 ;
    wire \LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_18 ;
    wire \LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_21 ;
    wire \LED_Blink_Inst.r_Count_5HZZ0Z_19 ;
    wire \LED_Blink_Inst.r_Count_5HZZ0Z_20 ;
    wire \LED_Blink_Inst.r_Count_5HZZ0Z_21 ;
    wire \LED_Blink_Inst.r_Count_5HZZ0Z_15 ;
    wire \LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_7 ;
    wire \LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_5 ;
    wire \LED_Blink_Inst.r_Count_5HZZ0Z_4 ;
    wire \LED_Blink_Inst.r_Count_5HZZ0Z_2 ;
    wire \LED_Blink_Inst.r_Count_5HZZ0Z_6 ;
    wire \LED_Blink_Inst.r_Count_5HZZ0Z_7 ;
    wire \LED_Blink_Inst.r_Count_5HZZ0Z_1 ;
    wire \LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_8 ;
    wire \LED_Blink_Inst.r_Count_5HZZ0Z_8 ;
    wire o_LED_2_c;
    wire \LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_13 ;
    wire \LED_Blink_Inst.r_Count_5HZZ0Z_13 ;
    wire \LED_Blink_Inst.r_Count_5HZZ0Z_18 ;
    wire \LED_Blink_Inst.r_Count_5HZZ0Z_5 ;
    wire \LED_Blink_Inst.r_Count_5HZZ0Z_3 ;
    wire \LED_Blink_Inst.un1_r_count_5hz_13_cascade_ ;
    wire \LED_Blink_Inst.un1_r_count_5hz_3 ;
    wire \LED_Blink_Inst.un1_r_count_5hz_11 ;
    wire \LED_Blink_Inst.r_Count_5HZZ0Z_11 ;
    wire \LED_Blink_Inst.un1_r_count_5hz_17_cascade_ ;
    wire \LED_Blink_Inst.r_Count_5HZZ0Z_0 ;
    wire \LED_Blink_Inst.un1_r_count_5hz_19_cascade_ ;
    wire \LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_17 ;
    wire \LED_Blink_Inst.r_Count_5HZZ0Z_17 ;
    wire \LED_Blink_Inst.r_Count_5HZZ0Z_9 ;
    wire \LED_Blink_Inst.r_Count_5HZZ0Z_14 ;
    wire \LED_Blink_Inst.r_Count_5HZZ0Z_16 ;
    wire \LED_Blink_Inst.r_Count_5HZZ0Z_12 ;
    wire \LED_Blink_Inst.un1_r_count_5hz_15 ;
    wire \LED_Blink_Inst.un1_r_count_5hz_19 ;
    wire \LED_Blink_Inst.un1_r_count_5hz_14 ;
    wire \LED_Blink_Inst.un1_r_count_5hz_15_cascade_ ;
    wire \LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_10 ;
    wire \LED_Blink_Inst.r_Count_5HZZ0Z_10 ;
    wire bfn_8_7_0_;
    wire \LED_Blink_Inst.un4_r_count_1hz_cry_1 ;
    wire \LED_Blink_Inst.un4_r_count_1hz_cry_2 ;
    wire \LED_Blink_Inst.un4_r_count_1hz_cry_3 ;
    wire \LED_Blink_Inst.un4_r_count_1hz_cry_4 ;
    wire \LED_Blink_Inst.un4_r_count_1hz_cry_5 ;
    wire \LED_Blink_Inst.un4_r_count_1hz_cry_6 ;
    wire \LED_Blink_Inst.un4_r_count_1hz_cry_7 ;
    wire \LED_Blink_Inst.un4_r_count_1hz_cry_8 ;
    wire bfn_8_8_0_;
    wire \LED_Blink_Inst.un4_r_count_1hz_cry_9 ;
    wire \LED_Blink_Inst.un4_r_count_1hz_cry_10 ;
    wire \LED_Blink_Inst.un4_r_count_1hz_cry_11 ;
    wire \LED_Blink_Inst.un4_r_count_1hz_cry_12 ;
    wire \LED_Blink_Inst.un4_r_count_1hz_cry_13 ;
    wire \LED_Blink_Inst.un4_r_count_1hz_cry_14 ;
    wire \LED_Blink_Inst.un4_r_count_1hz_cry_15 ;
    wire \LED_Blink_Inst.un4_r_count_1hz_cry_16 ;
    wire bfn_8_9_0_;
    wire \LED_Blink_Inst.un4_r_count_1hz_cry_17 ;
    wire \LED_Blink_Inst.un4_r_count_1hz_cry_18 ;
    wire \LED_Blink_Inst.un4_r_count_1hz_cry_19 ;
    wire \LED_Blink_Inst.un4_r_count_1hz_cry_20 ;
    wire \LED_Blink_Inst.un4_r_count_1hz_cry_21 ;
    wire \LED_Blink_Inst.un4_r_count_1hz_cry_22 ;
    wire \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_23_cascade_ ;
    wire \LED_Blink_Inst.r_Count_1HZZ0Z_13 ;
    wire \LED_Blink_Inst.r_Count_1HZZ0Z_10 ;
    wire \LED_Blink_Inst.r_Count_1HZZ0Z_15 ;
    wire \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_8 ;
    wire o_LED_4_c;
    wire \LED_Blink_Inst.r_Count_1HZZ0Z_5 ;
    wire \LED_Blink_Inst.r_Count_1HZZ0Z_6 ;
    wire \LED_Blink_Inst.r_Count_1HZZ0Z_7 ;
    wire \LED_Blink_Inst.r_Count_1HZZ0Z_4 ;
    wire \LED_Blink_Inst.r_Count_1HZZ0Z_0 ;
    wire \LED_Blink_Inst.r_Count_1HZZ0Z_3 ;
    wire \LED_Blink_Inst.r_Count_1HZZ0Z_2 ;
    wire \LED_Blink_Inst.r_Count_1HZZ0Z_8 ;
    wire \LED_Blink_Inst.r_Count_1HZZ0Z_1 ;
    wire \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_11 ;
    wire \LED_Blink_Inst.r_Count_1HZZ0Z_11 ;
    wire \LED_Blink_Inst.un1_r_count_1hz_13 ;
    wire \LED_Blink_Inst.un1_r_count_1hz_14_cascade_ ;
    wire \LED_Blink_Inst.un1_r_count_1hz_12 ;
    wire \LED_Blink_Inst.un1_r_count_1hz_21_cascade_ ;
    wire \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_12 ;
    wire \LED_Blink_Inst.r_Count_1HZZ0Z_12 ;
    wire \LED_Blink_Inst.r_Count_1HZZ0Z_22 ;
    wire \LED_Blink_Inst.r_Count_1HZZ0Z_19 ;
    wire \LED_Blink_Inst.r_Count_1HZZ0Z_23 ;
    wire \LED_Blink_Inst.r_Count_1HZZ0Z_14 ;
    wire \LED_Blink_Inst.un1_r_count_1hz_16_cascade_ ;
    wire \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_16 ;
    wire \LED_Blink_Inst.r_Count_1HZZ0Z_16 ;
    wire \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_9 ;
    wire \LED_Blink_Inst.r_Count_1HZZ0Z_9 ;
    wire \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_20 ;
    wire \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_18 ;
    wire \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_21 ;
    wire \LED_Blink_Inst.un1_r_count_1hz_21 ;
    wire \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_17 ;
    wire \LED_Blink_Inst.un1_r_count_1hz_17 ;
    wire \LED_Blink_Inst.un1_r_count_1hz_16 ;
    wire \LED_Blink_Inst.r_Count_1HZZ0Z_20 ;
    wire \LED_Blink_Inst.r_Count_1HZZ0Z_18 ;
    wire \LED_Blink_Inst.r_Count_1HZZ0Z_21 ;
    wire \LED_Blink_Inst.r_Count_1HZZ0Z_17 ;
    wire \LED_Blink_Inst.un1_r_count_1hz_15 ;
    wire bfn_11_3_0_;
    wire \LED_Blink_Inst.un6_r_count_10hz_cry_1 ;
    wire \LED_Blink_Inst.un6_r_count_10hz_cry_2 ;
    wire \LED_Blink_Inst.un6_r_count_10hz_cry_3 ;
    wire \LED_Blink_Inst.un6_r_count_10hz_cry_4 ;
    wire \LED_Blink_Inst.un6_r_count_10hz_cry_5 ;
    wire \LED_Blink_Inst.un6_r_count_10hz_cry_6 ;
    wire \LED_Blink_Inst.un6_r_count_10hz_cry_7 ;
    wire \LED_Blink_Inst.un6_r_count_10hz_cry_8 ;
    wire bfn_11_4_0_;
    wire \LED_Blink_Inst.un6_r_count_10hz_cry_9 ;
    wire \LED_Blink_Inst.un6_r_count_10hz_cry_10 ;
    wire \LED_Blink_Inst.un6_r_count_10hz_cry_11 ;
    wire \LED_Blink_Inst.un6_r_count_10hz_cry_12 ;
    wire \LED_Blink_Inst.un6_r_count_10hz_cry_13 ;
    wire \LED_Blink_Inst.un6_r_count_10hz_cry_14 ;
    wire \LED_Blink_Inst.un6_r_count_10hz_cry_15 ;
    wire \LED_Blink_Inst.un6_r_count_10hz_cry_16 ;
    wire bfn_11_5_0_;
    wire \LED_Blink_Inst.un6_r_count_10hz_cry_17 ;
    wire \LED_Blink_Inst.un6_r_count_10hz_cry_18 ;
    wire \LED_Blink_Inst.un6_r_count_10hz_cry_19 ;
    wire \LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_20_cascade_ ;
    wire \LED_Blink_Inst.r_Count_10HZZ0Z_20 ;
    wire \LED_Blink_Inst.r_Count_10HZZ0Z_19 ;
    wire \LED_Blink_Inst.r_Count_10HZZ0Z_18 ;
    wire \LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_17 ;
    wire \LED_Blink_Inst.r_Count_10HZZ0Z_17 ;
    wire \LED_Blink_Inst.un1_r_count_2hz_11 ;
    wire \LED_Blink_Inst.un1_r_count_2hz_12 ;
    wire \LED_Blink_Inst.un1_r_count_2hz_14_cascade_ ;
    wire \LED_Blink_Inst.un1_r_count_2hz_13 ;
    wire \LED_Blink_Inst.un1_r_count_2hz_20_cascade_ ;
    wire \LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_7 ;
    wire \LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_4 ;
    wire \LED_Blink_Inst.r_Count_10HZZ0Z_5 ;
    wire \LED_Blink_Inst.r_Count_10HZZ0Z_3 ;
    wire \LED_Blink_Inst.r_Count_10HZZ0Z_0 ;
    wire \LED_Blink_Inst.r_Count_10HZZ0Z_4 ;
    wire \LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_6 ;
    wire \LED_Blink_Inst.r_Count_10HZZ0Z_6 ;
    wire \LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_16 ;
    wire \LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_12 ;
    wire \LED_Blink_Inst.r_Count_10HZZ0Z_13 ;
    wire \LED_Blink_Inst.r_Count_10HZZ0Z_15 ;
    wire \LED_Blink_Inst.r_Count_10HZZ0Z_14 ;
    wire \LED_Blink_Inst.r_Count_10HZZ0Z_11 ;
    wire \LED_Blink_Inst.r_Count_10HZZ0Z_12 ;
    wire \LED_Blink_Inst.r_Count_10HZZ0Z_7 ;
    wire \LED_Blink_Inst.r_Count_10HZZ0Z_16 ;
    wire \LED_Blink_Inst.r_Count_10HZZ0Z_2 ;
    wire \LED_Blink_Inst.r_Count_10HZZ0Z_1 ;
    wire \LED_Blink_Inst.un1_r_count_10hz_12_cascade_ ;
    wire \LED_Blink_Inst.un1_r_count_10hz_2 ;
    wire \LED_Blink_Inst.r_Count_10HZZ0Z_8 ;
    wire \LED_Blink_Inst.r_Count_10HZZ0Z_10 ;
    wire \LED_Blink_Inst.un1_r_count_10hz_16_cascade_ ;
    wire \LED_Blink_Inst.un1_r_count_10hz_10 ;
    wire \LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_9 ;
    wire \LED_Blink_Inst.un1_r_count_10hz_18_cascade_ ;
    wire \LED_Blink_Inst.r_Count_10HZZ0Z_9 ;
    wire \LED_Blink_Inst.un1_r_count_10hz_14 ;
    wire \LED_Blink_Inst.un1_r_count_10hz_13 ;
    wire \LED_Blink_Inst.un1_r_count_10hz_18 ;
    wire o_LED_1_c;
    wire \LED_Blink_Inst.r_Count_2HZZ0Z_1 ;
    wire \LED_Blink_Inst.r_Count_2HZZ0Z_0 ;
    wire bfn_12_6_0_;
    wire \LED_Blink_Inst.r_Count_2HZZ0Z_2 ;
    wire \LED_Blink_Inst.un4_r_count_2hz_cry_1 ;
    wire \LED_Blink_Inst.r_Count_2HZZ0Z_3 ;
    wire \LED_Blink_Inst.un4_r_count_2hz_cry_2 ;
    wire \LED_Blink_Inst.r_Count_2HZZ0Z_4 ;
    wire \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_4 ;
    wire \LED_Blink_Inst.un4_r_count_2hz_cry_3 ;
    wire \LED_Blink_Inst.r_Count_2HZZ0Z_5 ;
    wire \LED_Blink_Inst.un4_r_count_2hz_cry_4 ;
    wire \LED_Blink_Inst.r_Count_2HZZ0Z_6 ;
    wire \LED_Blink_Inst.un4_r_count_2hz_cry_5 ;
    wire \LED_Blink_Inst.r_Count_2HZZ0Z_7 ;
    wire \LED_Blink_Inst.un4_r_count_2hz_cry_6 ;
    wire \LED_Blink_Inst.un4_r_count_2hz_cry_7 ;
    wire \LED_Blink_Inst.un4_r_count_2hz_cry_8 ;
    wire \LED_Blink_Inst.r_Count_2HZZ0Z_9 ;
    wire \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_9 ;
    wire bfn_12_7_0_;
    wire \LED_Blink_Inst.r_Count_2HZZ0Z_10 ;
    wire \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_10 ;
    wire \LED_Blink_Inst.un4_r_count_2hz_cry_9 ;
    wire \LED_Blink_Inst.r_Count_2HZZ0Z_11 ;
    wire \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_11 ;
    wire \LED_Blink_Inst.un4_r_count_2hz_cry_10 ;
    wire \LED_Blink_Inst.r_Count_2HZZ0Z_12 ;
    wire \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_12 ;
    wire \LED_Blink_Inst.un4_r_count_2hz_cry_11 ;
    wire \LED_Blink_Inst.un4_r_count_2hz_cry_12 ;
    wire \LED_Blink_Inst.r_Count_2HZZ0Z_14 ;
    wire \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_14 ;
    wire \LED_Blink_Inst.un4_r_count_2hz_cry_13 ;
    wire \LED_Blink_Inst.un4_r_count_2hz_cry_14 ;
    wire \LED_Blink_Inst.r_Count_2HZZ0Z_16 ;
    wire \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_16 ;
    wire \LED_Blink_Inst.un4_r_count_2hz_cry_15 ;
    wire \LED_Blink_Inst.un4_r_count_2hz_cry_16 ;
    wire bfn_12_8_0_;
    wire \LED_Blink_Inst.un4_r_count_2hz_cry_17 ;
    wire \LED_Blink_Inst.r_Count_2HZZ0Z_19 ;
    wire \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_19 ;
    wire \LED_Blink_Inst.un4_r_count_2hz_cry_18 ;
    wire \LED_Blink_Inst.r_Count_2HZZ0Z_20 ;
    wire \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_20 ;
    wire \LED_Blink_Inst.un4_r_count_2hz_cry_19 ;
    wire \LED_Blink_Inst.un4_r_count_2hz_cry_20 ;
    wire \LED_Blink_Inst.un4_r_count_2hz_cry_21 ;
    wire \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_22_cascade_ ;
    wire \LED_Blink_Inst.r_Count_2HZZ0Z_22 ;
    wire \LED_Blink_Inst.r_Count_2HZZ0Z_15 ;
    wire \LED_Blink_Inst.r_Count_2HZZ0Z_13 ;
    wire \LED_Blink_Inst.r_Count_2HZZ0Z_21 ;
    wire \LED_Blink_Inst.r_Count_2HZZ0Z_8 ;
    wire \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_17 ;
    wire \LED_Blink_Inst.r_Count_2HZZ0Z_17 ;
    wire \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_18 ;
    wire \LED_Blink_Inst.r_Count_2HZZ0Z_18 ;
    wire \LED_Blink_Inst.un1_r_count_2hz_15 ;
    wire \LED_Blink_Inst.un1_r_count_2hz_16 ;
    wire \LED_Blink_Inst.un1_r_count_2hz_20 ;
    wire o_LED_3_c;
    wire i_Clk_c_g;
    wire _gnd_net_;

    PRE_IO_GBUF i_Clk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__4821),
            .GLOBALBUFFEROUTPUT(i_Clk_c_g));
    IO_PAD i_Clk_ibuf_gb_io_iopad (
            .OE(N__4823),
            .DIN(N__4822),
            .DOUT(N__4821),
            .PACKAGEPIN(i_Clk));
    defparam i_Clk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam i_Clk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO i_Clk_ibuf_gb_io_preio (
            .PADOEN(N__4823),
            .PADOUT(N__4822),
            .PADIN(N__4821),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_LED_1_obuf_iopad (
            .OE(N__4812),
            .DIN(N__4811),
            .DOUT(N__4810),
            .PACKAGEPIN(o_LED_1));
    defparam o_LED_1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_LED_1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_LED_1_obuf_preio (
            .PADOEN(N__4812),
            .PADOUT(N__4811),
            .PADIN(N__4810),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3796),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_LED_2_obuf_iopad (
            .OE(N__4803),
            .DIN(N__4802),
            .DOUT(N__4801),
            .PACKAGEPIN(o_LED_2));
    defparam o_LED_2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_LED_2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_LED_2_obuf_preio (
            .PADOEN(N__4803),
            .PADOUT(N__4802),
            .PADIN(N__4801),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2360),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_LED_3_obuf_iopad (
            .OE(N__4794),
            .DIN(N__4793),
            .DOUT(N__4792),
            .PACKAGEPIN(o_LED_3));
    defparam o_LED_3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_LED_3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_LED_3_obuf_preio (
            .PADOEN(N__4794),
            .PADOUT(N__4793),
            .PADIN(N__4792),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4466),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_LED_4_obuf_iopad (
            .OE(N__4785),
            .DIN(N__4784),
            .DOUT(N__4783),
            .PACKAGEPIN(o_LED_4));
    defparam o_LED_4_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_LED_4_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_LED_4_obuf_preio (
            .PADOEN(N__4785),
            .PADOUT(N__4784),
            .PADIN(N__4783),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2933),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__1055 (
            .O(N__4766),
            .I(\LED_Blink_Inst.un4_r_count_2hz_cry_20 ));
    InMux I__1054 (
            .O(N__4763),
            .I(\LED_Blink_Inst.un4_r_count_2hz_cry_21 ));
    CascadeMux I__1053 (
            .O(N__4760),
            .I(\LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_22_cascade_ ));
    CascadeMux I__1052 (
            .O(N__4757),
            .I(N__4753));
    InMux I__1051 (
            .O(N__4756),
            .I(N__4750));
    InMux I__1050 (
            .O(N__4753),
            .I(N__4747));
    LocalMux I__1049 (
            .O(N__4750),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_22 ));
    LocalMux I__1048 (
            .O(N__4747),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_22 ));
    InMux I__1047 (
            .O(N__4742),
            .I(N__4738));
    InMux I__1046 (
            .O(N__4741),
            .I(N__4735));
    LocalMux I__1045 (
            .O(N__4738),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_15 ));
    LocalMux I__1044 (
            .O(N__4735),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_15 ));
    InMux I__1043 (
            .O(N__4730),
            .I(N__4726));
    InMux I__1042 (
            .O(N__4729),
            .I(N__4723));
    LocalMux I__1041 (
            .O(N__4726),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_13 ));
    LocalMux I__1040 (
            .O(N__4723),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_13 ));
    CascadeMux I__1039 (
            .O(N__4718),
            .I(N__4715));
    InMux I__1038 (
            .O(N__4715),
            .I(N__4709));
    InMux I__1037 (
            .O(N__4714),
            .I(N__4709));
    LocalMux I__1036 (
            .O(N__4709),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_21 ));
    InMux I__1035 (
            .O(N__4706),
            .I(N__4703));
    LocalMux I__1034 (
            .O(N__4703),
            .I(N__4699));
    InMux I__1033 (
            .O(N__4702),
            .I(N__4696));
    Odrv4 I__1032 (
            .O(N__4699),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_8 ));
    LocalMux I__1031 (
            .O(N__4696),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_8 ));
    CascadeMux I__1030 (
            .O(N__4691),
            .I(N__4688));
    InMux I__1029 (
            .O(N__4688),
            .I(N__4685));
    LocalMux I__1028 (
            .O(N__4685),
            .I(\LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_17 ));
    CascadeMux I__1027 (
            .O(N__4682),
            .I(N__4679));
    InMux I__1026 (
            .O(N__4679),
            .I(N__4675));
    InMux I__1025 (
            .O(N__4678),
            .I(N__4672));
    LocalMux I__1024 (
            .O(N__4675),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_17 ));
    LocalMux I__1023 (
            .O(N__4672),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_17 ));
    InMux I__1022 (
            .O(N__4667),
            .I(N__4664));
    LocalMux I__1021 (
            .O(N__4664),
            .I(\LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_18 ));
    InMux I__1020 (
            .O(N__4661),
            .I(N__4657));
    InMux I__1019 (
            .O(N__4660),
            .I(N__4654));
    LocalMux I__1018 (
            .O(N__4657),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_18 ));
    LocalMux I__1017 (
            .O(N__4654),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_18 ));
    InMux I__1016 (
            .O(N__4649),
            .I(N__4629));
    InMux I__1015 (
            .O(N__4648),
            .I(N__4629));
    InMux I__1014 (
            .O(N__4647),
            .I(N__4629));
    InMux I__1013 (
            .O(N__4646),
            .I(N__4626));
    InMux I__1012 (
            .O(N__4645),
            .I(N__4617));
    InMux I__1011 (
            .O(N__4644),
            .I(N__4617));
    InMux I__1010 (
            .O(N__4643),
            .I(N__4617));
    InMux I__1009 (
            .O(N__4642),
            .I(N__4617));
    InMux I__1008 (
            .O(N__4641),
            .I(N__4614));
    InMux I__1007 (
            .O(N__4640),
            .I(N__4603));
    InMux I__1006 (
            .O(N__4639),
            .I(N__4603));
    InMux I__1005 (
            .O(N__4638),
            .I(N__4603));
    InMux I__1004 (
            .O(N__4637),
            .I(N__4603));
    InMux I__1003 (
            .O(N__4636),
            .I(N__4603));
    LocalMux I__1002 (
            .O(N__4629),
            .I(\LED_Blink_Inst.un1_r_count_2hz_15 ));
    LocalMux I__1001 (
            .O(N__4626),
            .I(\LED_Blink_Inst.un1_r_count_2hz_15 ));
    LocalMux I__1000 (
            .O(N__4617),
            .I(\LED_Blink_Inst.un1_r_count_2hz_15 ));
    LocalMux I__999 (
            .O(N__4614),
            .I(\LED_Blink_Inst.un1_r_count_2hz_15 ));
    LocalMux I__998 (
            .O(N__4603),
            .I(\LED_Blink_Inst.un1_r_count_2hz_15 ));
    CascadeMux I__997 (
            .O(N__4592),
            .I(N__4587));
    CascadeMux I__996 (
            .O(N__4591),
            .I(N__4581));
    CascadeMux I__995 (
            .O(N__4590),
            .I(N__4575));
    InMux I__994 (
            .O(N__4587),
            .I(N__4563));
    InMux I__993 (
            .O(N__4586),
            .I(N__4563));
    InMux I__992 (
            .O(N__4585),
            .I(N__4563));
    InMux I__991 (
            .O(N__4584),
            .I(N__4552));
    InMux I__990 (
            .O(N__4581),
            .I(N__4552));
    InMux I__989 (
            .O(N__4580),
            .I(N__4552));
    InMux I__988 (
            .O(N__4579),
            .I(N__4552));
    InMux I__987 (
            .O(N__4578),
            .I(N__4552));
    InMux I__986 (
            .O(N__4575),
            .I(N__4541));
    InMux I__985 (
            .O(N__4574),
            .I(N__4541));
    InMux I__984 (
            .O(N__4573),
            .I(N__4541));
    InMux I__983 (
            .O(N__4572),
            .I(N__4541));
    InMux I__982 (
            .O(N__4571),
            .I(N__4541));
    InMux I__981 (
            .O(N__4570),
            .I(N__4538));
    LocalMux I__980 (
            .O(N__4563),
            .I(\LED_Blink_Inst.un1_r_count_2hz_16 ));
    LocalMux I__979 (
            .O(N__4552),
            .I(\LED_Blink_Inst.un1_r_count_2hz_16 ));
    LocalMux I__978 (
            .O(N__4541),
            .I(\LED_Blink_Inst.un1_r_count_2hz_16 ));
    LocalMux I__977 (
            .O(N__4538),
            .I(\LED_Blink_Inst.un1_r_count_2hz_16 ));
    CascadeMux I__976 (
            .O(N__4529),
            .I(N__4525));
    CascadeMux I__975 (
            .O(N__4528),
            .I(N__4521));
    InMux I__974 (
            .O(N__4525),
            .I(N__4506));
    InMux I__973 (
            .O(N__4524),
            .I(N__4506));
    InMux I__972 (
            .O(N__4521),
            .I(N__4499));
    InMux I__971 (
            .O(N__4520),
            .I(N__4499));
    InMux I__970 (
            .O(N__4519),
            .I(N__4499));
    InMux I__969 (
            .O(N__4518),
            .I(N__4496));
    InMux I__968 (
            .O(N__4517),
            .I(N__4489));
    InMux I__967 (
            .O(N__4516),
            .I(N__4489));
    InMux I__966 (
            .O(N__4515),
            .I(N__4489));
    InMux I__965 (
            .O(N__4514),
            .I(N__4480));
    InMux I__964 (
            .O(N__4513),
            .I(N__4480));
    InMux I__963 (
            .O(N__4512),
            .I(N__4480));
    InMux I__962 (
            .O(N__4511),
            .I(N__4480));
    LocalMux I__961 (
            .O(N__4506),
            .I(N__4475));
    LocalMux I__960 (
            .O(N__4499),
            .I(N__4475));
    LocalMux I__959 (
            .O(N__4496),
            .I(\LED_Blink_Inst.un1_r_count_2hz_20 ));
    LocalMux I__958 (
            .O(N__4489),
            .I(\LED_Blink_Inst.un1_r_count_2hz_20 ));
    LocalMux I__957 (
            .O(N__4480),
            .I(\LED_Blink_Inst.un1_r_count_2hz_20 ));
    Odrv4 I__956 (
            .O(N__4475),
            .I(\LED_Blink_Inst.un1_r_count_2hz_20 ));
    IoInMux I__955 (
            .O(N__4466),
            .I(N__4463));
    LocalMux I__954 (
            .O(N__4463),
            .I(N__4459));
    CascadeMux I__953 (
            .O(N__4462),
            .I(N__4456));
    Span4Mux_s0_h I__952 (
            .O(N__4459),
            .I(N__4453));
    InMux I__951 (
            .O(N__4456),
            .I(N__4450));
    Odrv4 I__950 (
            .O(N__4453),
            .I(o_LED_3_c));
    LocalMux I__949 (
            .O(N__4450),
            .I(o_LED_3_c));
    ClkMux I__948 (
            .O(N__4445),
            .I(N__4373));
    ClkMux I__947 (
            .O(N__4444),
            .I(N__4373));
    ClkMux I__946 (
            .O(N__4443),
            .I(N__4373));
    ClkMux I__945 (
            .O(N__4442),
            .I(N__4373));
    ClkMux I__944 (
            .O(N__4441),
            .I(N__4373));
    ClkMux I__943 (
            .O(N__4440),
            .I(N__4373));
    ClkMux I__942 (
            .O(N__4439),
            .I(N__4373));
    ClkMux I__941 (
            .O(N__4438),
            .I(N__4373));
    ClkMux I__940 (
            .O(N__4437),
            .I(N__4373));
    ClkMux I__939 (
            .O(N__4436),
            .I(N__4373));
    ClkMux I__938 (
            .O(N__4435),
            .I(N__4373));
    ClkMux I__937 (
            .O(N__4434),
            .I(N__4373));
    ClkMux I__936 (
            .O(N__4433),
            .I(N__4373));
    ClkMux I__935 (
            .O(N__4432),
            .I(N__4373));
    ClkMux I__934 (
            .O(N__4431),
            .I(N__4373));
    ClkMux I__933 (
            .O(N__4430),
            .I(N__4373));
    ClkMux I__932 (
            .O(N__4429),
            .I(N__4373));
    ClkMux I__931 (
            .O(N__4428),
            .I(N__4373));
    ClkMux I__930 (
            .O(N__4427),
            .I(N__4373));
    ClkMux I__929 (
            .O(N__4426),
            .I(N__4373));
    ClkMux I__928 (
            .O(N__4425),
            .I(N__4373));
    ClkMux I__927 (
            .O(N__4424),
            .I(N__4373));
    ClkMux I__926 (
            .O(N__4423),
            .I(N__4373));
    ClkMux I__925 (
            .O(N__4422),
            .I(N__4373));
    GlobalMux I__924 (
            .O(N__4373),
            .I(N__4370));
    gio2CtrlBuf I__923 (
            .O(N__4370),
            .I(i_Clk_c_g));
    InMux I__922 (
            .O(N__4367),
            .I(N__4363));
    InMux I__921 (
            .O(N__4366),
            .I(N__4360));
    LocalMux I__920 (
            .O(N__4363),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_12 ));
    LocalMux I__919 (
            .O(N__4360),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_12 ));
    CascadeMux I__918 (
            .O(N__4355),
            .I(N__4352));
    InMux I__917 (
            .O(N__4352),
            .I(N__4349));
    LocalMux I__916 (
            .O(N__4349),
            .I(N__4346));
    Span4Mux_v I__915 (
            .O(N__4346),
            .I(N__4343));
    Odrv4 I__914 (
            .O(N__4343),
            .I(\LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_12 ));
    InMux I__913 (
            .O(N__4340),
            .I(\LED_Blink_Inst.un4_r_count_2hz_cry_11 ));
    InMux I__912 (
            .O(N__4337),
            .I(\LED_Blink_Inst.un4_r_count_2hz_cry_12 ));
    InMux I__911 (
            .O(N__4334),
            .I(N__4330));
    InMux I__910 (
            .O(N__4333),
            .I(N__4327));
    LocalMux I__909 (
            .O(N__4330),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_14 ));
    LocalMux I__908 (
            .O(N__4327),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_14 ));
    InMux I__907 (
            .O(N__4322),
            .I(N__4319));
    LocalMux I__906 (
            .O(N__4319),
            .I(\LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_14 ));
    InMux I__905 (
            .O(N__4316),
            .I(\LED_Blink_Inst.un4_r_count_2hz_cry_13 ));
    InMux I__904 (
            .O(N__4313),
            .I(\LED_Blink_Inst.un4_r_count_2hz_cry_14 ));
    InMux I__903 (
            .O(N__4310),
            .I(N__4306));
    InMux I__902 (
            .O(N__4309),
            .I(N__4303));
    LocalMux I__901 (
            .O(N__4306),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_16 ));
    LocalMux I__900 (
            .O(N__4303),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_16 ));
    CascadeMux I__899 (
            .O(N__4298),
            .I(N__4295));
    InMux I__898 (
            .O(N__4295),
            .I(N__4292));
    LocalMux I__897 (
            .O(N__4292),
            .I(N__4289));
    Odrv4 I__896 (
            .O(N__4289),
            .I(\LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_16 ));
    InMux I__895 (
            .O(N__4286),
            .I(\LED_Blink_Inst.un4_r_count_2hz_cry_15 ));
    InMux I__894 (
            .O(N__4283),
            .I(bfn_12_8_0_));
    InMux I__893 (
            .O(N__4280),
            .I(\LED_Blink_Inst.un4_r_count_2hz_cry_17 ));
    InMux I__892 (
            .O(N__4277),
            .I(N__4273));
    InMux I__891 (
            .O(N__4276),
            .I(N__4270));
    LocalMux I__890 (
            .O(N__4273),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_19 ));
    LocalMux I__889 (
            .O(N__4270),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_19 ));
    CascadeMux I__888 (
            .O(N__4265),
            .I(N__4262));
    InMux I__887 (
            .O(N__4262),
            .I(N__4259));
    LocalMux I__886 (
            .O(N__4259),
            .I(\LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_19 ));
    InMux I__885 (
            .O(N__4256),
            .I(\LED_Blink_Inst.un4_r_count_2hz_cry_18 ));
    InMux I__884 (
            .O(N__4253),
            .I(N__4249));
    InMux I__883 (
            .O(N__4252),
            .I(N__4246));
    LocalMux I__882 (
            .O(N__4249),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_20 ));
    LocalMux I__881 (
            .O(N__4246),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_20 ));
    InMux I__880 (
            .O(N__4241),
            .I(N__4238));
    LocalMux I__879 (
            .O(N__4238),
            .I(\LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_20 ));
    InMux I__878 (
            .O(N__4235),
            .I(\LED_Blink_Inst.un4_r_count_2hz_cry_19 ));
    InMux I__877 (
            .O(N__4232),
            .I(N__4228));
    InMux I__876 (
            .O(N__4231),
            .I(N__4225));
    LocalMux I__875 (
            .O(N__4228),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_4 ));
    LocalMux I__874 (
            .O(N__4225),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_4 ));
    CascadeMux I__873 (
            .O(N__4220),
            .I(N__4217));
    InMux I__872 (
            .O(N__4217),
            .I(N__4214));
    LocalMux I__871 (
            .O(N__4214),
            .I(\LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_4 ));
    InMux I__870 (
            .O(N__4211),
            .I(\LED_Blink_Inst.un4_r_count_2hz_cry_3 ));
    CascadeMux I__869 (
            .O(N__4208),
            .I(N__4205));
    InMux I__868 (
            .O(N__4205),
            .I(N__4201));
    InMux I__867 (
            .O(N__4204),
            .I(N__4198));
    LocalMux I__866 (
            .O(N__4201),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_5 ));
    LocalMux I__865 (
            .O(N__4198),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_5 ));
    InMux I__864 (
            .O(N__4193),
            .I(\LED_Blink_Inst.un4_r_count_2hz_cry_4 ));
    InMux I__863 (
            .O(N__4190),
            .I(N__4186));
    InMux I__862 (
            .O(N__4189),
            .I(N__4183));
    LocalMux I__861 (
            .O(N__4186),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_6 ));
    LocalMux I__860 (
            .O(N__4183),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_6 ));
    InMux I__859 (
            .O(N__4178),
            .I(\LED_Blink_Inst.un4_r_count_2hz_cry_5 ));
    InMux I__858 (
            .O(N__4175),
            .I(N__4171));
    InMux I__857 (
            .O(N__4174),
            .I(N__4168));
    LocalMux I__856 (
            .O(N__4171),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_7 ));
    LocalMux I__855 (
            .O(N__4168),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_7 ));
    InMux I__854 (
            .O(N__4163),
            .I(\LED_Blink_Inst.un4_r_count_2hz_cry_6 ));
    InMux I__853 (
            .O(N__4160),
            .I(\LED_Blink_Inst.un4_r_count_2hz_cry_7 ));
    InMux I__852 (
            .O(N__4157),
            .I(N__4153));
    InMux I__851 (
            .O(N__4156),
            .I(N__4150));
    LocalMux I__850 (
            .O(N__4153),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_9 ));
    LocalMux I__849 (
            .O(N__4150),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_9 ));
    InMux I__848 (
            .O(N__4145),
            .I(N__4142));
    LocalMux I__847 (
            .O(N__4142),
            .I(\LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_9 ));
    InMux I__846 (
            .O(N__4139),
            .I(bfn_12_7_0_));
    InMux I__845 (
            .O(N__4136),
            .I(N__4132));
    InMux I__844 (
            .O(N__4135),
            .I(N__4129));
    LocalMux I__843 (
            .O(N__4132),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_10 ));
    LocalMux I__842 (
            .O(N__4129),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_10 ));
    CascadeMux I__841 (
            .O(N__4124),
            .I(N__4121));
    InMux I__840 (
            .O(N__4121),
            .I(N__4118));
    LocalMux I__839 (
            .O(N__4118),
            .I(\LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_10 ));
    InMux I__838 (
            .O(N__4115),
            .I(\LED_Blink_Inst.un4_r_count_2hz_cry_9 ));
    CascadeMux I__837 (
            .O(N__4112),
            .I(N__4109));
    InMux I__836 (
            .O(N__4109),
            .I(N__4105));
    InMux I__835 (
            .O(N__4108),
            .I(N__4102));
    LocalMux I__834 (
            .O(N__4105),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_11 ));
    LocalMux I__833 (
            .O(N__4102),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_11 ));
    InMux I__832 (
            .O(N__4097),
            .I(N__4094));
    LocalMux I__831 (
            .O(N__4094),
            .I(N__4091));
    Odrv4 I__830 (
            .O(N__4091),
            .I(\LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_11 ));
    InMux I__829 (
            .O(N__4088),
            .I(\LED_Blink_Inst.un4_r_count_2hz_cry_10 ));
    InMux I__828 (
            .O(N__4085),
            .I(N__4081));
    InMux I__827 (
            .O(N__4084),
            .I(N__4078));
    LocalMux I__826 (
            .O(N__4081),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_12 ));
    LocalMux I__825 (
            .O(N__4078),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_12 ));
    CascadeMux I__824 (
            .O(N__4073),
            .I(N__4069));
    InMux I__823 (
            .O(N__4072),
            .I(N__4066));
    InMux I__822 (
            .O(N__4069),
            .I(N__4063));
    LocalMux I__821 (
            .O(N__4066),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_7 ));
    LocalMux I__820 (
            .O(N__4063),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_7 ));
    InMux I__819 (
            .O(N__4058),
            .I(N__4054));
    InMux I__818 (
            .O(N__4057),
            .I(N__4051));
    LocalMux I__817 (
            .O(N__4054),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_16 ));
    LocalMux I__816 (
            .O(N__4051),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_16 ));
    InMux I__815 (
            .O(N__4046),
            .I(N__4042));
    InMux I__814 (
            .O(N__4045),
            .I(N__4039));
    LocalMux I__813 (
            .O(N__4042),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_2 ));
    LocalMux I__812 (
            .O(N__4039),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_2 ));
    InMux I__811 (
            .O(N__4034),
            .I(N__4029));
    InMux I__810 (
            .O(N__4033),
            .I(N__4026));
    InMux I__809 (
            .O(N__4032),
            .I(N__4023));
    LocalMux I__808 (
            .O(N__4029),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_1 ));
    LocalMux I__807 (
            .O(N__4026),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_1 ));
    LocalMux I__806 (
            .O(N__4023),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_1 ));
    CascadeMux I__805 (
            .O(N__4016),
            .I(\LED_Blink_Inst.un1_r_count_10hz_12_cascade_ ));
    InMux I__804 (
            .O(N__4013),
            .I(N__4010));
    LocalMux I__803 (
            .O(N__4010),
            .I(\LED_Blink_Inst.un1_r_count_10hz_2 ));
    InMux I__802 (
            .O(N__4007),
            .I(N__4003));
    InMux I__801 (
            .O(N__4006),
            .I(N__4000));
    LocalMux I__800 (
            .O(N__4003),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_8 ));
    LocalMux I__799 (
            .O(N__4000),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_8 ));
    InMux I__798 (
            .O(N__3995),
            .I(N__3991));
    InMux I__797 (
            .O(N__3994),
            .I(N__3988));
    LocalMux I__796 (
            .O(N__3991),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_10 ));
    LocalMux I__795 (
            .O(N__3988),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_10 ));
    CascadeMux I__794 (
            .O(N__3983),
            .I(\LED_Blink_Inst.un1_r_count_10hz_16_cascade_ ));
    InMux I__793 (
            .O(N__3980),
            .I(N__3977));
    LocalMux I__792 (
            .O(N__3977),
            .I(N__3974));
    Odrv4 I__791 (
            .O(N__3974),
            .I(\LED_Blink_Inst.un1_r_count_10hz_10 ));
    InMux I__790 (
            .O(N__3971),
            .I(N__3968));
    LocalMux I__789 (
            .O(N__3968),
            .I(\LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_9 ));
    CascadeMux I__788 (
            .O(N__3965),
            .I(\LED_Blink_Inst.un1_r_count_10hz_18_cascade_ ));
    InMux I__787 (
            .O(N__3962),
            .I(N__3958));
    InMux I__786 (
            .O(N__3961),
            .I(N__3955));
    LocalMux I__785 (
            .O(N__3958),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_9 ));
    LocalMux I__784 (
            .O(N__3955),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_9 ));
    CascadeMux I__783 (
            .O(N__3950),
            .I(N__3942));
    CascadeMux I__782 (
            .O(N__3949),
            .I(N__3936));
    CascadeMux I__781 (
            .O(N__3948),
            .I(N__3933));
    CascadeMux I__780 (
            .O(N__3947),
            .I(N__3929));
    CascadeMux I__779 (
            .O(N__3946),
            .I(N__3926));
    InMux I__778 (
            .O(N__3945),
            .I(N__3921));
    InMux I__777 (
            .O(N__3942),
            .I(N__3921));
    InMux I__776 (
            .O(N__3941),
            .I(N__3918));
    InMux I__775 (
            .O(N__3940),
            .I(N__3909));
    InMux I__774 (
            .O(N__3939),
            .I(N__3909));
    InMux I__773 (
            .O(N__3936),
            .I(N__3909));
    InMux I__772 (
            .O(N__3933),
            .I(N__3909));
    InMux I__771 (
            .O(N__3932),
            .I(N__3902));
    InMux I__770 (
            .O(N__3929),
            .I(N__3902));
    InMux I__769 (
            .O(N__3926),
            .I(N__3902));
    LocalMux I__768 (
            .O(N__3921),
            .I(\LED_Blink_Inst.un1_r_count_10hz_14 ));
    LocalMux I__767 (
            .O(N__3918),
            .I(\LED_Blink_Inst.un1_r_count_10hz_14 ));
    LocalMux I__766 (
            .O(N__3909),
            .I(\LED_Blink_Inst.un1_r_count_10hz_14 ));
    LocalMux I__765 (
            .O(N__3902),
            .I(\LED_Blink_Inst.un1_r_count_10hz_14 ));
    CascadeMux I__764 (
            .O(N__3893),
            .I(N__3889));
    CascadeMux I__763 (
            .O(N__3892),
            .I(N__3886));
    InMux I__762 (
            .O(N__3889),
            .I(N__3871));
    InMux I__761 (
            .O(N__3886),
            .I(N__3871));
    InMux I__760 (
            .O(N__3885),
            .I(N__3871));
    InMux I__759 (
            .O(N__3884),
            .I(N__3868));
    InMux I__758 (
            .O(N__3883),
            .I(N__3865));
    InMux I__757 (
            .O(N__3882),
            .I(N__3862));
    InMux I__756 (
            .O(N__3881),
            .I(N__3857));
    InMux I__755 (
            .O(N__3880),
            .I(N__3857));
    InMux I__754 (
            .O(N__3879),
            .I(N__3852));
    InMux I__753 (
            .O(N__3878),
            .I(N__3852));
    LocalMux I__752 (
            .O(N__3871),
            .I(N__3847));
    LocalMux I__751 (
            .O(N__3868),
            .I(N__3847));
    LocalMux I__750 (
            .O(N__3865),
            .I(\LED_Blink_Inst.un1_r_count_10hz_13 ));
    LocalMux I__749 (
            .O(N__3862),
            .I(\LED_Blink_Inst.un1_r_count_10hz_13 ));
    LocalMux I__748 (
            .O(N__3857),
            .I(\LED_Blink_Inst.un1_r_count_10hz_13 ));
    LocalMux I__747 (
            .O(N__3852),
            .I(\LED_Blink_Inst.un1_r_count_10hz_13 ));
    Odrv4 I__746 (
            .O(N__3847),
            .I(\LED_Blink_Inst.un1_r_count_10hz_13 ));
    InMux I__745 (
            .O(N__3836),
            .I(N__3825));
    InMux I__744 (
            .O(N__3835),
            .I(N__3820));
    InMux I__743 (
            .O(N__3834),
            .I(N__3820));
    InMux I__742 (
            .O(N__3833),
            .I(N__3815));
    InMux I__741 (
            .O(N__3832),
            .I(N__3815));
    InMux I__740 (
            .O(N__3831),
            .I(N__3806));
    InMux I__739 (
            .O(N__3830),
            .I(N__3806));
    InMux I__738 (
            .O(N__3829),
            .I(N__3806));
    InMux I__737 (
            .O(N__3828),
            .I(N__3806));
    LocalMux I__736 (
            .O(N__3825),
            .I(\LED_Blink_Inst.un1_r_count_10hz_18 ));
    LocalMux I__735 (
            .O(N__3820),
            .I(\LED_Blink_Inst.un1_r_count_10hz_18 ));
    LocalMux I__734 (
            .O(N__3815),
            .I(\LED_Blink_Inst.un1_r_count_10hz_18 ));
    LocalMux I__733 (
            .O(N__3806),
            .I(\LED_Blink_Inst.un1_r_count_10hz_18 ));
    CascadeMux I__732 (
            .O(N__3797),
            .I(N__3793));
    IoInMux I__731 (
            .O(N__3796),
            .I(N__3790));
    InMux I__730 (
            .O(N__3793),
            .I(N__3787));
    LocalMux I__729 (
            .O(N__3790),
            .I(o_LED_1_c));
    LocalMux I__728 (
            .O(N__3787),
            .I(o_LED_1_c));
    InMux I__727 (
            .O(N__3782),
            .I(N__3777));
    InMux I__726 (
            .O(N__3781),
            .I(N__3774));
    InMux I__725 (
            .O(N__3780),
            .I(N__3771));
    LocalMux I__724 (
            .O(N__3777),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_1 ));
    LocalMux I__723 (
            .O(N__3774),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_1 ));
    LocalMux I__722 (
            .O(N__3771),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_1 ));
    CascadeMux I__721 (
            .O(N__3764),
            .I(N__3758));
    InMux I__720 (
            .O(N__3763),
            .I(N__3755));
    InMux I__719 (
            .O(N__3762),
            .I(N__3750));
    InMux I__718 (
            .O(N__3761),
            .I(N__3750));
    InMux I__717 (
            .O(N__3758),
            .I(N__3747));
    LocalMux I__716 (
            .O(N__3755),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_0 ));
    LocalMux I__715 (
            .O(N__3750),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_0 ));
    LocalMux I__714 (
            .O(N__3747),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_0 ));
    InMux I__713 (
            .O(N__3740),
            .I(N__3736));
    InMux I__712 (
            .O(N__3739),
            .I(N__3733));
    LocalMux I__711 (
            .O(N__3736),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_2 ));
    LocalMux I__710 (
            .O(N__3733),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_2 ));
    InMux I__709 (
            .O(N__3728),
            .I(\LED_Blink_Inst.un4_r_count_2hz_cry_1 ));
    InMux I__708 (
            .O(N__3725),
            .I(N__3721));
    InMux I__707 (
            .O(N__3724),
            .I(N__3718));
    LocalMux I__706 (
            .O(N__3721),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_3 ));
    LocalMux I__705 (
            .O(N__3718),
            .I(\LED_Blink_Inst.r_Count_2HZZ0Z_3 ));
    InMux I__704 (
            .O(N__3713),
            .I(\LED_Blink_Inst.un4_r_count_2hz_cry_2 ));
    InMux I__703 (
            .O(N__3710),
            .I(N__3707));
    LocalMux I__702 (
            .O(N__3707),
            .I(\LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_4 ));
    InMux I__701 (
            .O(N__3704),
            .I(N__3700));
    InMux I__700 (
            .O(N__3703),
            .I(N__3697));
    LocalMux I__699 (
            .O(N__3700),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_5 ));
    LocalMux I__698 (
            .O(N__3697),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_5 ));
    InMux I__697 (
            .O(N__3692),
            .I(N__3688));
    InMux I__696 (
            .O(N__3691),
            .I(N__3685));
    LocalMux I__695 (
            .O(N__3688),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_3 ));
    LocalMux I__694 (
            .O(N__3685),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_3 ));
    CascadeMux I__693 (
            .O(N__3680),
            .I(N__3674));
    InMux I__692 (
            .O(N__3679),
            .I(N__3667));
    InMux I__691 (
            .O(N__3678),
            .I(N__3667));
    InMux I__690 (
            .O(N__3677),
            .I(N__3667));
    InMux I__689 (
            .O(N__3674),
            .I(N__3664));
    LocalMux I__688 (
            .O(N__3667),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_0 ));
    LocalMux I__687 (
            .O(N__3664),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_0 ));
    InMux I__686 (
            .O(N__3659),
            .I(N__3655));
    InMux I__685 (
            .O(N__3658),
            .I(N__3652));
    LocalMux I__684 (
            .O(N__3655),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_4 ));
    LocalMux I__683 (
            .O(N__3652),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_4 ));
    InMux I__682 (
            .O(N__3647),
            .I(N__3644));
    LocalMux I__681 (
            .O(N__3644),
            .I(\LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_6 ));
    InMux I__680 (
            .O(N__3641),
            .I(N__3637));
    InMux I__679 (
            .O(N__3640),
            .I(N__3634));
    LocalMux I__678 (
            .O(N__3637),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_6 ));
    LocalMux I__677 (
            .O(N__3634),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_6 ));
    InMux I__676 (
            .O(N__3629),
            .I(N__3626));
    LocalMux I__675 (
            .O(N__3626),
            .I(\LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_16 ));
    InMux I__674 (
            .O(N__3623),
            .I(N__3620));
    LocalMux I__673 (
            .O(N__3620),
            .I(\LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_12 ));
    InMux I__672 (
            .O(N__3617),
            .I(N__3613));
    InMux I__671 (
            .O(N__3616),
            .I(N__3610));
    LocalMux I__670 (
            .O(N__3613),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_13 ));
    LocalMux I__669 (
            .O(N__3610),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_13 ));
    InMux I__668 (
            .O(N__3605),
            .I(N__3601));
    InMux I__667 (
            .O(N__3604),
            .I(N__3598));
    LocalMux I__666 (
            .O(N__3601),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_15 ));
    LocalMux I__665 (
            .O(N__3598),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_15 ));
    CascadeMux I__664 (
            .O(N__3593),
            .I(N__3590));
    InMux I__663 (
            .O(N__3590),
            .I(N__3586));
    InMux I__662 (
            .O(N__3589),
            .I(N__3583));
    LocalMux I__661 (
            .O(N__3586),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_14 ));
    LocalMux I__660 (
            .O(N__3583),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_14 ));
    InMux I__659 (
            .O(N__3578),
            .I(N__3574));
    InMux I__658 (
            .O(N__3577),
            .I(N__3571));
    LocalMux I__657 (
            .O(N__3574),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_11 ));
    LocalMux I__656 (
            .O(N__3571),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_11 ));
    InMux I__655 (
            .O(N__3566),
            .I(N__3563));
    LocalMux I__654 (
            .O(N__3563),
            .I(\LED_Blink_Inst.un1_r_count_2hz_11 ));
    InMux I__653 (
            .O(N__3560),
            .I(N__3557));
    LocalMux I__652 (
            .O(N__3557),
            .I(\LED_Blink_Inst.un1_r_count_2hz_12 ));
    CascadeMux I__651 (
            .O(N__3554),
            .I(\LED_Blink_Inst.un1_r_count_2hz_14_cascade_ ));
    InMux I__650 (
            .O(N__3551),
            .I(N__3548));
    LocalMux I__649 (
            .O(N__3548),
            .I(\LED_Blink_Inst.un1_r_count_2hz_13 ));
    CascadeMux I__648 (
            .O(N__3545),
            .I(\LED_Blink_Inst.un1_r_count_2hz_20_cascade_ ));
    InMux I__647 (
            .O(N__3542),
            .I(N__3539));
    LocalMux I__646 (
            .O(N__3539),
            .I(\LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_7 ));
    InMux I__645 (
            .O(N__3536),
            .I(N__3533));
    LocalMux I__644 (
            .O(N__3533),
            .I(\LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_17 ));
    InMux I__643 (
            .O(N__3530),
            .I(N__3524));
    InMux I__642 (
            .O(N__3529),
            .I(N__3524));
    LocalMux I__641 (
            .O(N__3524),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_17 ));
    InMux I__640 (
            .O(N__3521),
            .I(\LED_Blink_Inst.un6_r_count_10hz_cry_13 ));
    InMux I__639 (
            .O(N__3518),
            .I(\LED_Blink_Inst.un6_r_count_10hz_cry_14 ));
    InMux I__638 (
            .O(N__3515),
            .I(\LED_Blink_Inst.un6_r_count_10hz_cry_15 ));
    InMux I__637 (
            .O(N__3512),
            .I(bfn_11_5_0_));
    InMux I__636 (
            .O(N__3509),
            .I(\LED_Blink_Inst.un6_r_count_10hz_cry_17 ));
    InMux I__635 (
            .O(N__3506),
            .I(\LED_Blink_Inst.un6_r_count_10hz_cry_18 ));
    InMux I__634 (
            .O(N__3503),
            .I(\LED_Blink_Inst.un6_r_count_10hz_cry_19 ));
    CascadeMux I__633 (
            .O(N__3500),
            .I(\LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_20_cascade_ ));
    InMux I__632 (
            .O(N__3497),
            .I(N__3491));
    InMux I__631 (
            .O(N__3496),
            .I(N__3491));
    LocalMux I__630 (
            .O(N__3491),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_20 ));
    CascadeMux I__629 (
            .O(N__3488),
            .I(N__3485));
    InMux I__628 (
            .O(N__3485),
            .I(N__3479));
    InMux I__627 (
            .O(N__3484),
            .I(N__3479));
    LocalMux I__626 (
            .O(N__3479),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_19 ));
    InMux I__625 (
            .O(N__3476),
            .I(N__3470));
    InMux I__624 (
            .O(N__3475),
            .I(N__3470));
    LocalMux I__623 (
            .O(N__3470),
            .I(\LED_Blink_Inst.r_Count_10HZZ0Z_18 ));
    InMux I__622 (
            .O(N__3467),
            .I(\LED_Blink_Inst.un6_r_count_10hz_cry_4 ));
    InMux I__621 (
            .O(N__3464),
            .I(\LED_Blink_Inst.un6_r_count_10hz_cry_5 ));
    InMux I__620 (
            .O(N__3461),
            .I(\LED_Blink_Inst.un6_r_count_10hz_cry_6 ));
    InMux I__619 (
            .O(N__3458),
            .I(\LED_Blink_Inst.un6_r_count_10hz_cry_7 ));
    InMux I__618 (
            .O(N__3455),
            .I(bfn_11_4_0_));
    InMux I__617 (
            .O(N__3452),
            .I(\LED_Blink_Inst.un6_r_count_10hz_cry_9 ));
    InMux I__616 (
            .O(N__3449),
            .I(\LED_Blink_Inst.un6_r_count_10hz_cry_10 ));
    InMux I__615 (
            .O(N__3446),
            .I(\LED_Blink_Inst.un6_r_count_10hz_cry_11 ));
    InMux I__614 (
            .O(N__3443),
            .I(\LED_Blink_Inst.un6_r_count_10hz_cry_12 ));
    InMux I__613 (
            .O(N__3440),
            .I(N__3437));
    LocalMux I__612 (
            .O(N__3437),
            .I(\LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_18 ));
    InMux I__611 (
            .O(N__3434),
            .I(N__3431));
    LocalMux I__610 (
            .O(N__3431),
            .I(\LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_21 ));
    InMux I__609 (
            .O(N__3428),
            .I(N__3415));
    InMux I__608 (
            .O(N__3427),
            .I(N__3406));
    InMux I__607 (
            .O(N__3426),
            .I(N__3406));
    InMux I__606 (
            .O(N__3425),
            .I(N__3406));
    InMux I__605 (
            .O(N__3424),
            .I(N__3406));
    InMux I__604 (
            .O(N__3423),
            .I(N__3397));
    InMux I__603 (
            .O(N__3422),
            .I(N__3397));
    InMux I__602 (
            .O(N__3421),
            .I(N__3397));
    InMux I__601 (
            .O(N__3420),
            .I(N__3397));
    InMux I__600 (
            .O(N__3419),
            .I(N__3392));
    InMux I__599 (
            .O(N__3418),
            .I(N__3392));
    LocalMux I__598 (
            .O(N__3415),
            .I(\LED_Blink_Inst.un1_r_count_1hz_21 ));
    LocalMux I__597 (
            .O(N__3406),
            .I(\LED_Blink_Inst.un1_r_count_1hz_21 ));
    LocalMux I__596 (
            .O(N__3397),
            .I(\LED_Blink_Inst.un1_r_count_1hz_21 ));
    LocalMux I__595 (
            .O(N__3392),
            .I(\LED_Blink_Inst.un1_r_count_1hz_21 ));
    InMux I__594 (
            .O(N__3383),
            .I(N__3380));
    LocalMux I__593 (
            .O(N__3380),
            .I(\LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_17 ));
    CascadeMux I__592 (
            .O(N__3377),
            .I(N__3366));
    CascadeMux I__591 (
            .O(N__3376),
            .I(N__3363));
    CascadeMux I__590 (
            .O(N__3375),
            .I(N__3360));
    CascadeMux I__589 (
            .O(N__3374),
            .I(N__3357));
    CascadeMux I__588 (
            .O(N__3373),
            .I(N__3354));
    CascadeMux I__587 (
            .O(N__3372),
            .I(N__3351));
    InMux I__586 (
            .O(N__3371),
            .I(N__3347));
    CascadeMux I__585 (
            .O(N__3370),
            .I(N__3342));
    InMux I__584 (
            .O(N__3369),
            .I(N__3339));
    InMux I__583 (
            .O(N__3366),
            .I(N__3334));
    InMux I__582 (
            .O(N__3363),
            .I(N__3334));
    InMux I__581 (
            .O(N__3360),
            .I(N__3329));
    InMux I__580 (
            .O(N__3357),
            .I(N__3329));
    InMux I__579 (
            .O(N__3354),
            .I(N__3326));
    InMux I__578 (
            .O(N__3351),
            .I(N__3321));
    InMux I__577 (
            .O(N__3350),
            .I(N__3321));
    LocalMux I__576 (
            .O(N__3347),
            .I(N__3318));
    InMux I__575 (
            .O(N__3346),
            .I(N__3311));
    InMux I__574 (
            .O(N__3345),
            .I(N__3311));
    InMux I__573 (
            .O(N__3342),
            .I(N__3311));
    LocalMux I__572 (
            .O(N__3339),
            .I(N__3308));
    LocalMux I__571 (
            .O(N__3334),
            .I(N__3303));
    LocalMux I__570 (
            .O(N__3329),
            .I(N__3303));
    LocalMux I__569 (
            .O(N__3326),
            .I(N__3296));
    LocalMux I__568 (
            .O(N__3321),
            .I(N__3296));
    Span4Mux_h I__567 (
            .O(N__3318),
            .I(N__3296));
    LocalMux I__566 (
            .O(N__3311),
            .I(\LED_Blink_Inst.un1_r_count_1hz_17 ));
    Odrv4 I__565 (
            .O(N__3308),
            .I(\LED_Blink_Inst.un1_r_count_1hz_17 ));
    Odrv12 I__564 (
            .O(N__3303),
            .I(\LED_Blink_Inst.un1_r_count_1hz_17 ));
    Odrv4 I__563 (
            .O(N__3296),
            .I(\LED_Blink_Inst.un1_r_count_1hz_17 ));
    InMux I__562 (
            .O(N__3287),
            .I(N__3270));
    InMux I__561 (
            .O(N__3286),
            .I(N__3270));
    InMux I__560 (
            .O(N__3285),
            .I(N__3270));
    InMux I__559 (
            .O(N__3284),
            .I(N__3270));
    InMux I__558 (
            .O(N__3283),
            .I(N__3265));
    InMux I__557 (
            .O(N__3282),
            .I(N__3256));
    InMux I__556 (
            .O(N__3281),
            .I(N__3256));
    InMux I__555 (
            .O(N__3280),
            .I(N__3256));
    InMux I__554 (
            .O(N__3279),
            .I(N__3256));
    LocalMux I__553 (
            .O(N__3270),
            .I(N__3253));
    InMux I__552 (
            .O(N__3269),
            .I(N__3248));
    InMux I__551 (
            .O(N__3268),
            .I(N__3248));
    LocalMux I__550 (
            .O(N__3265),
            .I(\LED_Blink_Inst.un1_r_count_1hz_16 ));
    LocalMux I__549 (
            .O(N__3256),
            .I(\LED_Blink_Inst.un1_r_count_1hz_16 ));
    Odrv4 I__548 (
            .O(N__3253),
            .I(\LED_Blink_Inst.un1_r_count_1hz_16 ));
    LocalMux I__547 (
            .O(N__3248),
            .I(\LED_Blink_Inst.un1_r_count_1hz_16 ));
    InMux I__546 (
            .O(N__3239),
            .I(N__3235));
    InMux I__545 (
            .O(N__3238),
            .I(N__3232));
    LocalMux I__544 (
            .O(N__3235),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_20 ));
    LocalMux I__543 (
            .O(N__3232),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_20 ));
    InMux I__542 (
            .O(N__3227),
            .I(N__3223));
    InMux I__541 (
            .O(N__3226),
            .I(N__3220));
    LocalMux I__540 (
            .O(N__3223),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_18 ));
    LocalMux I__539 (
            .O(N__3220),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_18 ));
    CascadeMux I__538 (
            .O(N__3215),
            .I(N__3211));
    InMux I__537 (
            .O(N__3214),
            .I(N__3208));
    InMux I__536 (
            .O(N__3211),
            .I(N__3205));
    LocalMux I__535 (
            .O(N__3208),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_21 ));
    LocalMux I__534 (
            .O(N__3205),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_21 ));
    InMux I__533 (
            .O(N__3200),
            .I(N__3196));
    InMux I__532 (
            .O(N__3199),
            .I(N__3193));
    LocalMux I__531 (
            .O(N__3196),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_17 ));
    LocalMux I__530 (
            .O(N__3193),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_17 ));
    InMux I__529 (
            .O(N__3188),
            .I(N__3185));
    LocalMux I__528 (
            .O(N__3185),
            .I(\LED_Blink_Inst.un1_r_count_1hz_15 ));
    InMux I__527 (
            .O(N__3182),
            .I(\LED_Blink_Inst.un6_r_count_10hz_cry_1 ));
    InMux I__526 (
            .O(N__3179),
            .I(\LED_Blink_Inst.un6_r_count_10hz_cry_2 ));
    InMux I__525 (
            .O(N__3176),
            .I(\LED_Blink_Inst.un6_r_count_10hz_cry_3 ));
    InMux I__524 (
            .O(N__3173),
            .I(N__3166));
    InMux I__523 (
            .O(N__3172),
            .I(N__3166));
    InMux I__522 (
            .O(N__3171),
            .I(N__3163));
    LocalMux I__521 (
            .O(N__3166),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_1 ));
    LocalMux I__520 (
            .O(N__3163),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_1 ));
    CascadeMux I__519 (
            .O(N__3158),
            .I(N__3155));
    InMux I__518 (
            .O(N__3155),
            .I(N__3152));
    LocalMux I__517 (
            .O(N__3152),
            .I(\LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_11 ));
    InMux I__516 (
            .O(N__3149),
            .I(N__3145));
    InMux I__515 (
            .O(N__3148),
            .I(N__3142));
    LocalMux I__514 (
            .O(N__3145),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_11 ));
    LocalMux I__513 (
            .O(N__3142),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_11 ));
    InMux I__512 (
            .O(N__3137),
            .I(N__3134));
    LocalMux I__511 (
            .O(N__3134),
            .I(N__3131));
    Odrv4 I__510 (
            .O(N__3131),
            .I(\LED_Blink_Inst.un1_r_count_1hz_13 ));
    CascadeMux I__509 (
            .O(N__3128),
            .I(\LED_Blink_Inst.un1_r_count_1hz_14_cascade_ ));
    InMux I__508 (
            .O(N__3125),
            .I(N__3122));
    LocalMux I__507 (
            .O(N__3122),
            .I(\LED_Blink_Inst.un1_r_count_1hz_12 ));
    CascadeMux I__506 (
            .O(N__3119),
            .I(\LED_Blink_Inst.un1_r_count_1hz_21_cascade_ ));
    InMux I__505 (
            .O(N__3116),
            .I(N__3113));
    LocalMux I__504 (
            .O(N__3113),
            .I(\LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_12 ));
    InMux I__503 (
            .O(N__3110),
            .I(N__3106));
    InMux I__502 (
            .O(N__3109),
            .I(N__3103));
    LocalMux I__501 (
            .O(N__3106),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_12 ));
    LocalMux I__500 (
            .O(N__3103),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_12 ));
    InMux I__499 (
            .O(N__3098),
            .I(N__3094));
    InMux I__498 (
            .O(N__3097),
            .I(N__3091));
    LocalMux I__497 (
            .O(N__3094),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_22 ));
    LocalMux I__496 (
            .O(N__3091),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_22 ));
    InMux I__495 (
            .O(N__3086),
            .I(N__3082));
    InMux I__494 (
            .O(N__3085),
            .I(N__3079));
    LocalMux I__493 (
            .O(N__3082),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_19 ));
    LocalMux I__492 (
            .O(N__3079),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_19 ));
    CascadeMux I__491 (
            .O(N__3074),
            .I(N__3071));
    InMux I__490 (
            .O(N__3071),
            .I(N__3067));
    InMux I__489 (
            .O(N__3070),
            .I(N__3064));
    LocalMux I__488 (
            .O(N__3067),
            .I(N__3061));
    LocalMux I__487 (
            .O(N__3064),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_23 ));
    Odrv4 I__486 (
            .O(N__3061),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_23 ));
    InMux I__485 (
            .O(N__3056),
            .I(N__3052));
    InMux I__484 (
            .O(N__3055),
            .I(N__3049));
    LocalMux I__483 (
            .O(N__3052),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_14 ));
    LocalMux I__482 (
            .O(N__3049),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_14 ));
    CascadeMux I__481 (
            .O(N__3044),
            .I(\LED_Blink_Inst.un1_r_count_1hz_16_cascade_ ));
    InMux I__480 (
            .O(N__3041),
            .I(N__3038));
    LocalMux I__479 (
            .O(N__3038),
            .I(\LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_16 ));
    CascadeMux I__478 (
            .O(N__3035),
            .I(N__3032));
    InMux I__477 (
            .O(N__3032),
            .I(N__3028));
    InMux I__476 (
            .O(N__3031),
            .I(N__3025));
    LocalMux I__475 (
            .O(N__3028),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_16 ));
    LocalMux I__474 (
            .O(N__3025),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_16 ));
    InMux I__473 (
            .O(N__3020),
            .I(N__3017));
    LocalMux I__472 (
            .O(N__3017),
            .I(\LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_9 ));
    InMux I__471 (
            .O(N__3014),
            .I(N__3010));
    InMux I__470 (
            .O(N__3013),
            .I(N__3007));
    LocalMux I__469 (
            .O(N__3010),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_9 ));
    LocalMux I__468 (
            .O(N__3007),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_9 ));
    InMux I__467 (
            .O(N__3002),
            .I(N__2999));
    LocalMux I__466 (
            .O(N__2999),
            .I(\LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_20 ));
    InMux I__465 (
            .O(N__2996),
            .I(\LED_Blink_Inst.un4_r_count_1hz_cry_22 ));
    CascadeMux I__464 (
            .O(N__2993),
            .I(\LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_23_cascade_ ));
    InMux I__463 (
            .O(N__2990),
            .I(N__2987));
    LocalMux I__462 (
            .O(N__2987),
            .I(N__2983));
    InMux I__461 (
            .O(N__2986),
            .I(N__2980));
    Odrv4 I__460 (
            .O(N__2983),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_13 ));
    LocalMux I__459 (
            .O(N__2980),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_13 ));
    InMux I__458 (
            .O(N__2975),
            .I(N__2972));
    LocalMux I__457 (
            .O(N__2972),
            .I(N__2968));
    InMux I__456 (
            .O(N__2971),
            .I(N__2965));
    Odrv4 I__455 (
            .O(N__2968),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_10 ));
    LocalMux I__454 (
            .O(N__2965),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_10 ));
    CascadeMux I__453 (
            .O(N__2960),
            .I(N__2957));
    InMux I__452 (
            .O(N__2957),
            .I(N__2953));
    CascadeMux I__451 (
            .O(N__2956),
            .I(N__2950));
    LocalMux I__450 (
            .O(N__2953),
            .I(N__2947));
    InMux I__449 (
            .O(N__2950),
            .I(N__2944));
    Odrv4 I__448 (
            .O(N__2947),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_15 ));
    LocalMux I__447 (
            .O(N__2944),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_15 ));
    InMux I__446 (
            .O(N__2939),
            .I(N__2936));
    LocalMux I__445 (
            .O(N__2936),
            .I(\LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_8 ));
    IoInMux I__444 (
            .O(N__2933),
            .I(N__2930));
    LocalMux I__443 (
            .O(N__2930),
            .I(N__2926));
    CascadeMux I__442 (
            .O(N__2929),
            .I(N__2923));
    Span4Mux_s2_h I__441 (
            .O(N__2926),
            .I(N__2920));
    InMux I__440 (
            .O(N__2923),
            .I(N__2917));
    Odrv4 I__439 (
            .O(N__2920),
            .I(o_LED_4_c));
    LocalMux I__438 (
            .O(N__2917),
            .I(o_LED_4_c));
    InMux I__437 (
            .O(N__2912),
            .I(N__2908));
    InMux I__436 (
            .O(N__2911),
            .I(N__2905));
    LocalMux I__435 (
            .O(N__2908),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_5 ));
    LocalMux I__434 (
            .O(N__2905),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_5 ));
    InMux I__433 (
            .O(N__2900),
            .I(N__2896));
    InMux I__432 (
            .O(N__2899),
            .I(N__2893));
    LocalMux I__431 (
            .O(N__2896),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_6 ));
    LocalMux I__430 (
            .O(N__2893),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_6 ));
    CascadeMux I__429 (
            .O(N__2888),
            .I(N__2885));
    InMux I__428 (
            .O(N__2885),
            .I(N__2881));
    InMux I__427 (
            .O(N__2884),
            .I(N__2878));
    LocalMux I__426 (
            .O(N__2881),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_7 ));
    LocalMux I__425 (
            .O(N__2878),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_7 ));
    InMux I__424 (
            .O(N__2873),
            .I(N__2869));
    InMux I__423 (
            .O(N__2872),
            .I(N__2866));
    LocalMux I__422 (
            .O(N__2869),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_4 ));
    LocalMux I__421 (
            .O(N__2866),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_4 ));
    CascadeMux I__420 (
            .O(N__2861),
            .I(N__2857));
    CascadeMux I__419 (
            .O(N__2860),
            .I(N__2852));
    InMux I__418 (
            .O(N__2857),
            .I(N__2847));
    InMux I__417 (
            .O(N__2856),
            .I(N__2847));
    InMux I__416 (
            .O(N__2855),
            .I(N__2844));
    InMux I__415 (
            .O(N__2852),
            .I(N__2841));
    LocalMux I__414 (
            .O(N__2847),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_0 ));
    LocalMux I__413 (
            .O(N__2844),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_0 ));
    LocalMux I__412 (
            .O(N__2841),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_0 ));
    InMux I__411 (
            .O(N__2834),
            .I(N__2830));
    InMux I__410 (
            .O(N__2833),
            .I(N__2827));
    LocalMux I__409 (
            .O(N__2830),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_3 ));
    LocalMux I__408 (
            .O(N__2827),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_3 ));
    InMux I__407 (
            .O(N__2822),
            .I(N__2818));
    InMux I__406 (
            .O(N__2821),
            .I(N__2815));
    LocalMux I__405 (
            .O(N__2818),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_2 ));
    LocalMux I__404 (
            .O(N__2815),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_2 ));
    CascadeMux I__403 (
            .O(N__2810),
            .I(N__2807));
    InMux I__402 (
            .O(N__2807),
            .I(N__2803));
    InMux I__401 (
            .O(N__2806),
            .I(N__2800));
    LocalMux I__400 (
            .O(N__2803),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_8 ));
    LocalMux I__399 (
            .O(N__2800),
            .I(\LED_Blink_Inst.r_Count_1HZZ0Z_8 ));
    InMux I__398 (
            .O(N__2795),
            .I(\LED_Blink_Inst.un4_r_count_1hz_cry_13 ));
    InMux I__397 (
            .O(N__2792),
            .I(\LED_Blink_Inst.un4_r_count_1hz_cry_14 ));
    InMux I__396 (
            .O(N__2789),
            .I(\LED_Blink_Inst.un4_r_count_1hz_cry_15 ));
    InMux I__395 (
            .O(N__2786),
            .I(bfn_8_9_0_));
    InMux I__394 (
            .O(N__2783),
            .I(\LED_Blink_Inst.un4_r_count_1hz_cry_17 ));
    InMux I__393 (
            .O(N__2780),
            .I(\LED_Blink_Inst.un4_r_count_1hz_cry_18 ));
    InMux I__392 (
            .O(N__2777),
            .I(\LED_Blink_Inst.un4_r_count_1hz_cry_19 ));
    InMux I__391 (
            .O(N__2774),
            .I(\LED_Blink_Inst.un4_r_count_1hz_cry_20 ));
    InMux I__390 (
            .O(N__2771),
            .I(\LED_Blink_Inst.un4_r_count_1hz_cry_21 ));
    InMux I__389 (
            .O(N__2768),
            .I(\LED_Blink_Inst.un4_r_count_1hz_cry_4 ));
    InMux I__388 (
            .O(N__2765),
            .I(\LED_Blink_Inst.un4_r_count_1hz_cry_5 ));
    InMux I__387 (
            .O(N__2762),
            .I(\LED_Blink_Inst.un4_r_count_1hz_cry_6 ));
    InMux I__386 (
            .O(N__2759),
            .I(\LED_Blink_Inst.un4_r_count_1hz_cry_7 ));
    InMux I__385 (
            .O(N__2756),
            .I(bfn_8_8_0_));
    InMux I__384 (
            .O(N__2753),
            .I(\LED_Blink_Inst.un4_r_count_1hz_cry_9 ));
    InMux I__383 (
            .O(N__2750),
            .I(\LED_Blink_Inst.un4_r_count_1hz_cry_10 ));
    InMux I__382 (
            .O(N__2747),
            .I(\LED_Blink_Inst.un4_r_count_1hz_cry_11 ));
    InMux I__381 (
            .O(N__2744),
            .I(\LED_Blink_Inst.un4_r_count_1hz_cry_12 ));
    InMux I__380 (
            .O(N__2741),
            .I(N__2738));
    LocalMux I__379 (
            .O(N__2738),
            .I(\LED_Blink_Inst.un1_r_count_5hz_11 ));
    InMux I__378 (
            .O(N__2735),
            .I(N__2731));
    InMux I__377 (
            .O(N__2734),
            .I(N__2728));
    LocalMux I__376 (
            .O(N__2731),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_11 ));
    LocalMux I__375 (
            .O(N__2728),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_11 ));
    CascadeMux I__374 (
            .O(N__2723),
            .I(\LED_Blink_Inst.un1_r_count_5hz_17_cascade_ ));
    CascadeMux I__373 (
            .O(N__2720),
            .I(N__2714));
    InMux I__372 (
            .O(N__2719),
            .I(N__2711));
    InMux I__371 (
            .O(N__2718),
            .I(N__2706));
    InMux I__370 (
            .O(N__2717),
            .I(N__2706));
    InMux I__369 (
            .O(N__2714),
            .I(N__2703));
    LocalMux I__368 (
            .O(N__2711),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_0 ));
    LocalMux I__367 (
            .O(N__2706),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_0 ));
    LocalMux I__366 (
            .O(N__2703),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_0 ));
    CascadeMux I__365 (
            .O(N__2696),
            .I(\LED_Blink_Inst.un1_r_count_5hz_19_cascade_ ));
    InMux I__364 (
            .O(N__2693),
            .I(N__2690));
    LocalMux I__363 (
            .O(N__2690),
            .I(\LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_17 ));
    CascadeMux I__362 (
            .O(N__2687),
            .I(N__2684));
    InMux I__361 (
            .O(N__2684),
            .I(N__2680));
    InMux I__360 (
            .O(N__2683),
            .I(N__2677));
    LocalMux I__359 (
            .O(N__2680),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_17 ));
    LocalMux I__358 (
            .O(N__2677),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_17 ));
    InMux I__357 (
            .O(N__2672),
            .I(N__2668));
    InMux I__356 (
            .O(N__2671),
            .I(N__2665));
    LocalMux I__355 (
            .O(N__2668),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_9 ));
    LocalMux I__354 (
            .O(N__2665),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_9 ));
    InMux I__353 (
            .O(N__2660),
            .I(N__2656));
    InMux I__352 (
            .O(N__2659),
            .I(N__2653));
    LocalMux I__351 (
            .O(N__2656),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_14 ));
    LocalMux I__350 (
            .O(N__2653),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_14 ));
    CascadeMux I__349 (
            .O(N__2648),
            .I(N__2645));
    InMux I__348 (
            .O(N__2645),
            .I(N__2641));
    InMux I__347 (
            .O(N__2644),
            .I(N__2638));
    LocalMux I__346 (
            .O(N__2641),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_16 ));
    LocalMux I__345 (
            .O(N__2638),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_16 ));
    InMux I__344 (
            .O(N__2633),
            .I(N__2629));
    InMux I__343 (
            .O(N__2632),
            .I(N__2626));
    LocalMux I__342 (
            .O(N__2629),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_12 ));
    LocalMux I__341 (
            .O(N__2626),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_12 ));
    CascadeMux I__340 (
            .O(N__2621),
            .I(N__2613));
    InMux I__339 (
            .O(N__2620),
            .I(N__2609));
    CascadeMux I__338 (
            .O(N__2619),
            .I(N__2606));
    InMux I__337 (
            .O(N__2618),
            .I(N__2597));
    InMux I__336 (
            .O(N__2617),
            .I(N__2597));
    InMux I__335 (
            .O(N__2616),
            .I(N__2597));
    InMux I__334 (
            .O(N__2613),
            .I(N__2597));
    CascadeMux I__333 (
            .O(N__2612),
            .I(N__2592));
    LocalMux I__332 (
            .O(N__2609),
            .I(N__2589));
    InMux I__331 (
            .O(N__2606),
            .I(N__2586));
    LocalMux I__330 (
            .O(N__2597),
            .I(N__2583));
    InMux I__329 (
            .O(N__2596),
            .I(N__2578));
    InMux I__328 (
            .O(N__2595),
            .I(N__2578));
    InMux I__327 (
            .O(N__2592),
            .I(N__2575));
    Odrv4 I__326 (
            .O(N__2589),
            .I(\LED_Blink_Inst.un1_r_count_5hz_15 ));
    LocalMux I__325 (
            .O(N__2586),
            .I(\LED_Blink_Inst.un1_r_count_5hz_15 ));
    Odrv4 I__324 (
            .O(N__2583),
            .I(\LED_Blink_Inst.un1_r_count_5hz_15 ));
    LocalMux I__323 (
            .O(N__2578),
            .I(\LED_Blink_Inst.un1_r_count_5hz_15 ));
    LocalMux I__322 (
            .O(N__2575),
            .I(\LED_Blink_Inst.un1_r_count_5hz_15 ));
    CascadeMux I__321 (
            .O(N__2564),
            .I(N__2557));
    CascadeMux I__320 (
            .O(N__2563),
            .I(N__2552));
    CascadeMux I__319 (
            .O(N__2562),
            .I(N__2549));
    CascadeMux I__318 (
            .O(N__2561),
            .I(N__2545));
    InMux I__317 (
            .O(N__2560),
            .I(N__2539));
    InMux I__316 (
            .O(N__2557),
            .I(N__2539));
    InMux I__315 (
            .O(N__2556),
            .I(N__2530));
    InMux I__314 (
            .O(N__2555),
            .I(N__2530));
    InMux I__313 (
            .O(N__2552),
            .I(N__2530));
    InMux I__312 (
            .O(N__2549),
            .I(N__2530));
    InMux I__311 (
            .O(N__2548),
            .I(N__2523));
    InMux I__310 (
            .O(N__2545),
            .I(N__2523));
    InMux I__309 (
            .O(N__2544),
            .I(N__2523));
    LocalMux I__308 (
            .O(N__2539),
            .I(\LED_Blink_Inst.un1_r_count_5hz_19 ));
    LocalMux I__307 (
            .O(N__2530),
            .I(\LED_Blink_Inst.un1_r_count_5hz_19 ));
    LocalMux I__306 (
            .O(N__2523),
            .I(\LED_Blink_Inst.un1_r_count_5hz_19 ));
    InMux I__305 (
            .O(N__2516),
            .I(N__2504));
    InMux I__304 (
            .O(N__2515),
            .I(N__2504));
    InMux I__303 (
            .O(N__2514),
            .I(N__2504));
    InMux I__302 (
            .O(N__2513),
            .I(N__2504));
    LocalMux I__301 (
            .O(N__2504),
            .I(N__2495));
    InMux I__300 (
            .O(N__2503),
            .I(N__2486));
    InMux I__299 (
            .O(N__2502),
            .I(N__2486));
    InMux I__298 (
            .O(N__2501),
            .I(N__2486));
    InMux I__297 (
            .O(N__2500),
            .I(N__2486));
    InMux I__296 (
            .O(N__2499),
            .I(N__2481));
    InMux I__295 (
            .O(N__2498),
            .I(N__2481));
    Odrv4 I__294 (
            .O(N__2495),
            .I(\LED_Blink_Inst.un1_r_count_5hz_14 ));
    LocalMux I__293 (
            .O(N__2486),
            .I(\LED_Blink_Inst.un1_r_count_5hz_14 ));
    LocalMux I__292 (
            .O(N__2481),
            .I(\LED_Blink_Inst.un1_r_count_5hz_14 ));
    CascadeMux I__291 (
            .O(N__2474),
            .I(\LED_Blink_Inst.un1_r_count_5hz_15_cascade_ ));
    InMux I__290 (
            .O(N__2471),
            .I(N__2468));
    LocalMux I__289 (
            .O(N__2468),
            .I(\LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_10 ));
    InMux I__288 (
            .O(N__2465),
            .I(N__2461));
    InMux I__287 (
            .O(N__2464),
            .I(N__2458));
    LocalMux I__286 (
            .O(N__2461),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_10 ));
    LocalMux I__285 (
            .O(N__2458),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_10 ));
    InMux I__284 (
            .O(N__2453),
            .I(\LED_Blink_Inst.un4_r_count_1hz_cry_1 ));
    InMux I__283 (
            .O(N__2450),
            .I(\LED_Blink_Inst.un4_r_count_1hz_cry_2 ));
    InMux I__282 (
            .O(N__2447),
            .I(\LED_Blink_Inst.un4_r_count_1hz_cry_3 ));
    InMux I__281 (
            .O(N__2444),
            .I(N__2440));
    InMux I__280 (
            .O(N__2443),
            .I(N__2437));
    LocalMux I__279 (
            .O(N__2440),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_4 ));
    LocalMux I__278 (
            .O(N__2437),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_4 ));
    InMux I__277 (
            .O(N__2432),
            .I(N__2428));
    InMux I__276 (
            .O(N__2431),
            .I(N__2425));
    LocalMux I__275 (
            .O(N__2428),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_2 ));
    LocalMux I__274 (
            .O(N__2425),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_2 ));
    CascadeMux I__273 (
            .O(N__2420),
            .I(N__2417));
    InMux I__272 (
            .O(N__2417),
            .I(N__2413));
    InMux I__271 (
            .O(N__2416),
            .I(N__2410));
    LocalMux I__270 (
            .O(N__2413),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_6 ));
    LocalMux I__269 (
            .O(N__2410),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_6 ));
    InMux I__268 (
            .O(N__2405),
            .I(N__2401));
    InMux I__267 (
            .O(N__2404),
            .I(N__2398));
    LocalMux I__266 (
            .O(N__2401),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_7 ));
    LocalMux I__265 (
            .O(N__2398),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_7 ));
    InMux I__264 (
            .O(N__2393),
            .I(N__2386));
    InMux I__263 (
            .O(N__2392),
            .I(N__2386));
    InMux I__262 (
            .O(N__2391),
            .I(N__2383));
    LocalMux I__261 (
            .O(N__2386),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_1 ));
    LocalMux I__260 (
            .O(N__2383),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_1 ));
    InMux I__259 (
            .O(N__2378),
            .I(N__2375));
    LocalMux I__258 (
            .O(N__2375),
            .I(\LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_8 ));
    InMux I__257 (
            .O(N__2372),
            .I(N__2368));
    InMux I__256 (
            .O(N__2371),
            .I(N__2365));
    LocalMux I__255 (
            .O(N__2368),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_8 ));
    LocalMux I__254 (
            .O(N__2365),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_8 ));
    IoInMux I__253 (
            .O(N__2360),
            .I(N__2357));
    LocalMux I__252 (
            .O(N__2357),
            .I(N__2353));
    CascadeMux I__251 (
            .O(N__2356),
            .I(N__2350));
    Span4Mux_s3_h I__250 (
            .O(N__2353),
            .I(N__2347));
    InMux I__249 (
            .O(N__2350),
            .I(N__2344));
    Odrv4 I__248 (
            .O(N__2347),
            .I(o_LED_2_c));
    LocalMux I__247 (
            .O(N__2344),
            .I(o_LED_2_c));
    InMux I__246 (
            .O(N__2339),
            .I(N__2336));
    LocalMux I__245 (
            .O(N__2336),
            .I(\LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_13 ));
    InMux I__244 (
            .O(N__2333),
            .I(N__2329));
    InMux I__243 (
            .O(N__2332),
            .I(N__2326));
    LocalMux I__242 (
            .O(N__2329),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_13 ));
    LocalMux I__241 (
            .O(N__2326),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_13 ));
    InMux I__240 (
            .O(N__2321),
            .I(N__2317));
    InMux I__239 (
            .O(N__2320),
            .I(N__2314));
    LocalMux I__238 (
            .O(N__2317),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_18 ));
    LocalMux I__237 (
            .O(N__2314),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_18 ));
    InMux I__236 (
            .O(N__2309),
            .I(N__2305));
    InMux I__235 (
            .O(N__2308),
            .I(N__2302));
    LocalMux I__234 (
            .O(N__2305),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_5 ));
    LocalMux I__233 (
            .O(N__2302),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_5 ));
    InMux I__232 (
            .O(N__2297),
            .I(N__2293));
    InMux I__231 (
            .O(N__2296),
            .I(N__2290));
    LocalMux I__230 (
            .O(N__2293),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_3 ));
    LocalMux I__229 (
            .O(N__2290),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_3 ));
    CascadeMux I__228 (
            .O(N__2285),
            .I(\LED_Blink_Inst.un1_r_count_5hz_13_cascade_ ));
    InMux I__227 (
            .O(N__2282),
            .I(N__2279));
    LocalMux I__226 (
            .O(N__2279),
            .I(\LED_Blink_Inst.un1_r_count_5hz_3 ));
    InMux I__225 (
            .O(N__2276),
            .I(\LED_Blink_Inst.un4_r_count_5hz_cry_17 ));
    InMux I__224 (
            .O(N__2273),
            .I(\LED_Blink_Inst.un4_r_count_5hz_cry_18 ));
    InMux I__223 (
            .O(N__2270),
            .I(\LED_Blink_Inst.un4_r_count_5hz_cry_19 ));
    InMux I__222 (
            .O(N__2267),
            .I(\LED_Blink_Inst.un4_r_count_5hz_cry_20 ));
    InMux I__221 (
            .O(N__2264),
            .I(N__2261));
    LocalMux I__220 (
            .O(N__2261),
            .I(\LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_18 ));
    InMux I__219 (
            .O(N__2258),
            .I(N__2255));
    LocalMux I__218 (
            .O(N__2255),
            .I(\LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_21 ));
    InMux I__217 (
            .O(N__2252),
            .I(N__2246));
    InMux I__216 (
            .O(N__2251),
            .I(N__2246));
    LocalMux I__215 (
            .O(N__2246),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_19 ));
    InMux I__214 (
            .O(N__2243),
            .I(N__2237));
    InMux I__213 (
            .O(N__2242),
            .I(N__2237));
    LocalMux I__212 (
            .O(N__2237),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_20 ));
    CascadeMux I__211 (
            .O(N__2234),
            .I(N__2230));
    InMux I__210 (
            .O(N__2233),
            .I(N__2225));
    InMux I__209 (
            .O(N__2230),
            .I(N__2225));
    LocalMux I__208 (
            .O(N__2225),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_21 ));
    InMux I__207 (
            .O(N__2222),
            .I(N__2218));
    InMux I__206 (
            .O(N__2221),
            .I(N__2215));
    LocalMux I__205 (
            .O(N__2218),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_15 ));
    LocalMux I__204 (
            .O(N__2215),
            .I(\LED_Blink_Inst.r_Count_5HZZ0Z_15 ));
    InMux I__203 (
            .O(N__2210),
            .I(N__2207));
    LocalMux I__202 (
            .O(N__2207),
            .I(\LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_7 ));
    InMux I__201 (
            .O(N__2204),
            .I(N__2201));
    LocalMux I__200 (
            .O(N__2201),
            .I(\LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_5 ));
    InMux I__199 (
            .O(N__2198),
            .I(bfn_7_6_0_));
    InMux I__198 (
            .O(N__2195),
            .I(\LED_Blink_Inst.un4_r_count_5hz_cry_9 ));
    InMux I__197 (
            .O(N__2192),
            .I(\LED_Blink_Inst.un4_r_count_5hz_cry_10 ));
    InMux I__196 (
            .O(N__2189),
            .I(\LED_Blink_Inst.un4_r_count_5hz_cry_11 ));
    InMux I__195 (
            .O(N__2186),
            .I(\LED_Blink_Inst.un4_r_count_5hz_cry_12 ));
    InMux I__194 (
            .O(N__2183),
            .I(\LED_Blink_Inst.un4_r_count_5hz_cry_13 ));
    InMux I__193 (
            .O(N__2180),
            .I(\LED_Blink_Inst.un4_r_count_5hz_cry_14 ));
    InMux I__192 (
            .O(N__2177),
            .I(\LED_Blink_Inst.un4_r_count_5hz_cry_15 ));
    InMux I__191 (
            .O(N__2174),
            .I(bfn_7_7_0_));
    InMux I__190 (
            .O(N__2171),
            .I(\LED_Blink_Inst.un4_r_count_5hz_cry_1 ));
    InMux I__189 (
            .O(N__2168),
            .I(\LED_Blink_Inst.un4_r_count_5hz_cry_2 ));
    InMux I__188 (
            .O(N__2165),
            .I(\LED_Blink_Inst.un4_r_count_5hz_cry_3 ));
    InMux I__187 (
            .O(N__2162),
            .I(\LED_Blink_Inst.un4_r_count_5hz_cry_4 ));
    InMux I__186 (
            .O(N__2159),
            .I(\LED_Blink_Inst.un4_r_count_5hz_cry_5 ));
    InMux I__185 (
            .O(N__2156),
            .I(\LED_Blink_Inst.un4_r_count_5hz_cry_6 ));
    InMux I__184 (
            .O(N__2153),
            .I(\LED_Blink_Inst.un4_r_count_5hz_cry_7 ));
    defparam IN_MUX_bfv_11_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_3_0_));
    defparam IN_MUX_bfv_11_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_4_0_ (
            .carryinitin(\LED_Blink_Inst.un6_r_count_10hz_cry_8 ),
            .carryinitout(bfn_11_4_0_));
    defparam IN_MUX_bfv_11_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_5_0_ (
            .carryinitin(\LED_Blink_Inst.un6_r_count_10hz_cry_16 ),
            .carryinitout(bfn_11_5_0_));
    defparam IN_MUX_bfv_7_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_5_0_));
    defparam IN_MUX_bfv_7_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_6_0_ (
            .carryinitin(\LED_Blink_Inst.un4_r_count_5hz_cry_8 ),
            .carryinitout(bfn_7_6_0_));
    defparam IN_MUX_bfv_7_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_7_0_ (
            .carryinitin(\LED_Blink_Inst.un4_r_count_5hz_cry_16 ),
            .carryinitout(bfn_7_7_0_));
    defparam IN_MUX_bfv_12_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_6_0_));
    defparam IN_MUX_bfv_12_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_7_0_ (
            .carryinitin(\LED_Blink_Inst.un4_r_count_2hz_cry_8 ),
            .carryinitout(bfn_12_7_0_));
    defparam IN_MUX_bfv_12_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_8_0_ (
            .carryinitin(\LED_Blink_Inst.un4_r_count_2hz_cry_16 ),
            .carryinitout(bfn_12_8_0_));
    defparam IN_MUX_bfv_8_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_7_0_));
    defparam IN_MUX_bfv_8_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_8_0_ (
            .carryinitin(\LED_Blink_Inst.un4_r_count_1hz_cry_8 ),
            .carryinitout(bfn_8_8_0_));
    defparam IN_MUX_bfv_8_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_9_0_ (
            .carryinitin(\LED_Blink_Inst.un4_r_count_1hz_cry_16 ),
            .carryinitout(bfn_8_9_0_));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \LED_Blink_Inst.un4_r_count_5hz_cry_1_c_LC_7_5_0 .C_ON=1'b1;
    defparam \LED_Blink_Inst.un4_r_count_5hz_cry_1_c_LC_7_5_0 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.un4_r_count_5hz_cry_1_c_LC_7_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \LED_Blink_Inst.un4_r_count_5hz_cry_1_c_LC_7_5_0  (
            .in0(_gnd_net_),
            .in1(N__2391),
            .in2(N__2720),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_5_0_),
            .carryout(\LED_Blink_Inst.un4_r_count_5hz_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_2_LC_7_5_1 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_5HZ_2_LC_7_5_1 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_5HZ_2_LC_7_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_2_LC_7_5_1  (
            .in0(_gnd_net_),
            .in1(N__2431),
            .in2(_gnd_net_),
            .in3(N__2171),
            .lcout(\LED_Blink_Inst.r_Count_5HZZ0Z_2 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_5hz_cry_1 ),
            .carryout(\LED_Blink_Inst.un4_r_count_5hz_cry_2 ),
            .clk(N__4428),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_3_LC_7_5_2 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_5HZ_3_LC_7_5_2 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_5HZ_3_LC_7_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_3_LC_7_5_2  (
            .in0(_gnd_net_),
            .in1(N__2296),
            .in2(_gnd_net_),
            .in3(N__2168),
            .lcout(\LED_Blink_Inst.r_Count_5HZZ0Z_3 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_5hz_cry_2 ),
            .carryout(\LED_Blink_Inst.un4_r_count_5hz_cry_3 ),
            .clk(N__4428),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_4_LC_7_5_3 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_5HZ_4_LC_7_5_3 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_5HZ_4_LC_7_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_4_LC_7_5_3  (
            .in0(_gnd_net_),
            .in1(N__2443),
            .in2(_gnd_net_),
            .in3(N__2165),
            .lcout(\LED_Blink_Inst.r_Count_5HZZ0Z_4 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_5hz_cry_3 ),
            .carryout(\LED_Blink_Inst.un4_r_count_5hz_cry_4 ),
            .clk(N__4428),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_RNO_0_5_LC_7_5_4 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_5HZ_RNO_0_5_LC_7_5_4 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_5HZ_RNO_0_5_LC_7_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_RNO_0_5_LC_7_5_4  (
            .in0(_gnd_net_),
            .in1(N__2308),
            .in2(_gnd_net_),
            .in3(N__2162),
            .lcout(\LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_5hz_cry_4 ),
            .carryout(\LED_Blink_Inst.un4_r_count_5hz_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_6_LC_7_5_5 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_5HZ_6_LC_7_5_5 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_5HZ_6_LC_7_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_6_LC_7_5_5  (
            .in0(_gnd_net_),
            .in1(N__2416),
            .in2(_gnd_net_),
            .in3(N__2159),
            .lcout(\LED_Blink_Inst.r_Count_5HZZ0Z_6 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_5hz_cry_5 ),
            .carryout(\LED_Blink_Inst.un4_r_count_5hz_cry_6 ),
            .clk(N__4428),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_RNO_0_7_LC_7_5_6 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_5HZ_RNO_0_7_LC_7_5_6 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_5HZ_RNO_0_7_LC_7_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_RNO_0_7_LC_7_5_6  (
            .in0(_gnd_net_),
            .in1(N__2404),
            .in2(_gnd_net_),
            .in3(N__2156),
            .lcout(\LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_5hz_cry_6 ),
            .carryout(\LED_Blink_Inst.un4_r_count_5hz_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_RNO_0_8_LC_7_5_7 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_5HZ_RNO_0_8_LC_7_5_7 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_5HZ_RNO_0_8_LC_7_5_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_RNO_0_8_LC_7_5_7  (
            .in0(_gnd_net_),
            .in1(N__2372),
            .in2(_gnd_net_),
            .in3(N__2153),
            .lcout(\LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_5hz_cry_7 ),
            .carryout(\LED_Blink_Inst.un4_r_count_5hz_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_9_LC_7_6_0 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_5HZ_9_LC_7_6_0 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_5HZ_9_LC_7_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_9_LC_7_6_0  (
            .in0(_gnd_net_),
            .in1(N__2671),
            .in2(_gnd_net_),
            .in3(N__2198),
            .lcout(\LED_Blink_Inst.r_Count_5HZZ0Z_9 ),
            .ltout(),
            .carryin(bfn_7_6_0_),
            .carryout(\LED_Blink_Inst.un4_r_count_5hz_cry_9 ),
            .clk(N__4425),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_RNO_0_10_LC_7_6_1 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_5HZ_RNO_0_10_LC_7_6_1 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_5HZ_RNO_0_10_LC_7_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_RNO_0_10_LC_7_6_1  (
            .in0(_gnd_net_),
            .in1(N__2464),
            .in2(_gnd_net_),
            .in3(N__2195),
            .lcout(\LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_5hz_cry_9 ),
            .carryout(\LED_Blink_Inst.un4_r_count_5hz_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_11_LC_7_6_2 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_5HZ_11_LC_7_6_2 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_5HZ_11_LC_7_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_11_LC_7_6_2  (
            .in0(_gnd_net_),
            .in1(N__2734),
            .in2(_gnd_net_),
            .in3(N__2192),
            .lcout(\LED_Blink_Inst.r_Count_5HZZ0Z_11 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_5hz_cry_10 ),
            .carryout(\LED_Blink_Inst.un4_r_count_5hz_cry_11 ),
            .clk(N__4425),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_12_LC_7_6_3 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_5HZ_12_LC_7_6_3 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_5HZ_12_LC_7_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_12_LC_7_6_3  (
            .in0(_gnd_net_),
            .in1(N__2632),
            .in2(_gnd_net_),
            .in3(N__2189),
            .lcout(\LED_Blink_Inst.r_Count_5HZZ0Z_12 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_5hz_cry_11 ),
            .carryout(\LED_Blink_Inst.un4_r_count_5hz_cry_12 ),
            .clk(N__4425),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_RNO_0_13_LC_7_6_4 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_5HZ_RNO_0_13_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_5HZ_RNO_0_13_LC_7_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_RNO_0_13_LC_7_6_4  (
            .in0(_gnd_net_),
            .in1(N__2332),
            .in2(_gnd_net_),
            .in3(N__2186),
            .lcout(\LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_5hz_cry_12 ),
            .carryout(\LED_Blink_Inst.un4_r_count_5hz_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_14_LC_7_6_5 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_5HZ_14_LC_7_6_5 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_5HZ_14_LC_7_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_14_LC_7_6_5  (
            .in0(_gnd_net_),
            .in1(N__2659),
            .in2(_gnd_net_),
            .in3(N__2183),
            .lcout(\LED_Blink_Inst.r_Count_5HZZ0Z_14 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_5hz_cry_13 ),
            .carryout(\LED_Blink_Inst.un4_r_count_5hz_cry_14 ),
            .clk(N__4425),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_15_LC_7_6_6 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_5HZ_15_LC_7_6_6 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_5HZ_15_LC_7_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_15_LC_7_6_6  (
            .in0(_gnd_net_),
            .in1(N__2221),
            .in2(_gnd_net_),
            .in3(N__2180),
            .lcout(\LED_Blink_Inst.r_Count_5HZZ0Z_15 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_5hz_cry_14 ),
            .carryout(\LED_Blink_Inst.un4_r_count_5hz_cry_15 ),
            .clk(N__4425),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_16_LC_7_6_7 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_5HZ_16_LC_7_6_7 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_5HZ_16_LC_7_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_16_LC_7_6_7  (
            .in0(_gnd_net_),
            .in1(N__2644),
            .in2(_gnd_net_),
            .in3(N__2177),
            .lcout(\LED_Blink_Inst.r_Count_5HZZ0Z_16 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_5hz_cry_15 ),
            .carryout(\LED_Blink_Inst.un4_r_count_5hz_cry_16 ),
            .clk(N__4425),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_RNO_0_17_LC_7_7_0 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_5HZ_RNO_0_17_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_5HZ_RNO_0_17_LC_7_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_RNO_0_17_LC_7_7_0  (
            .in0(_gnd_net_),
            .in1(N__2683),
            .in2(_gnd_net_),
            .in3(N__2174),
            .lcout(\LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(bfn_7_7_0_),
            .carryout(\LED_Blink_Inst.un4_r_count_5hz_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_RNO_0_18_LC_7_7_1 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_5HZ_RNO_0_18_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_5HZ_RNO_0_18_LC_7_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_RNO_0_18_LC_7_7_1  (
            .in0(_gnd_net_),
            .in1(N__2321),
            .in2(_gnd_net_),
            .in3(N__2276),
            .lcout(\LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_5hz_cry_17 ),
            .carryout(\LED_Blink_Inst.un4_r_count_5hz_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_19_LC_7_7_2 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_5HZ_19_LC_7_7_2 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_5HZ_19_LC_7_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_19_LC_7_7_2  (
            .in0(_gnd_net_),
            .in1(N__2251),
            .in2(_gnd_net_),
            .in3(N__2273),
            .lcout(\LED_Blink_Inst.r_Count_5HZZ0Z_19 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_5hz_cry_18 ),
            .carryout(\LED_Blink_Inst.un4_r_count_5hz_cry_19 ),
            .clk(N__4423),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_20_LC_7_7_3 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_5HZ_20_LC_7_7_3 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_5HZ_20_LC_7_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_20_LC_7_7_3  (
            .in0(_gnd_net_),
            .in1(N__2242),
            .in2(_gnd_net_),
            .in3(N__2270),
            .lcout(\LED_Blink_Inst.r_Count_5HZZ0Z_20 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_5hz_cry_19 ),
            .carryout(\LED_Blink_Inst.un4_r_count_5hz_cry_20 ),
            .clk(N__4423),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_RNO_0_21_LC_7_7_4 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_5HZ_RNO_0_21_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_5HZ_RNO_0_21_LC_7_7_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_RNO_0_21_LC_7_7_4  (
            .in0(_gnd_net_),
            .in1(N__2233),
            .in2(_gnd_net_),
            .in3(N__2267),
            .lcout(\LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_18_LC_7_7_5 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_5HZ_18_LC_7_7_5 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_5HZ_18_LC_7_7_5 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_18_LC_7_7_5  (
            .in0(N__2498),
            .in1(N__2264),
            .in2(N__2619),
            .in3(N__2560),
            .lcout(\LED_Blink_Inst.r_Count_5HZZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4423),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_21_LC_7_7_6 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_5HZ_21_LC_7_7_6 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_5HZ_21_LC_7_7_6 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_21_LC_7_7_6  (
            .in0(N__2620),
            .in1(N__2499),
            .in2(N__2564),
            .in3(N__2258),
            .lcout(\LED_Blink_Inst.r_Count_5HZZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4423),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_RNIH2F11_21_LC_7_7_7 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_5HZ_RNIH2F11_21_LC_7_7_7 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_5HZ_RNIH2F11_21_LC_7_7_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_RNIH2F11_21_LC_7_7_7  (
            .in0(N__2252),
            .in1(N__2243),
            .in2(N__2234),
            .in3(N__2222),
            .lcout(\LED_Blink_Inst.un1_r_count_5hz_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_7_LC_8_5_0 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_5HZ_7_LC_8_5_0 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_5HZ_7_LC_8_5_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_7_LC_8_5_0  (
            .in0(N__2514),
            .in1(N__2616),
            .in2(N__2562),
            .in3(N__2210),
            .lcout(\LED_Blink_Inst.r_Count_5HZZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4433),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_5_LC_8_5_1 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_5HZ_5_LC_8_5_1 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_5HZ_5_LC_8_5_1 .LUT_INIT=16'b0010101010101010;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_5_LC_8_5_1  (
            .in0(N__2204),
            .in1(N__2513),
            .in2(N__2621),
            .in3(N__2555),
            .lcout(\LED_Blink_Inst.r_Count_5HZZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4433),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_RNI96LC_1_LC_8_5_2 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_5HZ_RNI96LC_1_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_5HZ_RNI96LC_1_LC_8_5_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_RNI96LC_1_LC_8_5_2  (
            .in0(N__2444),
            .in1(N__2432),
            .in2(N__2420),
            .in3(N__2392),
            .lcout(\LED_Blink_Inst.un1_r_count_5hz_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_RNITRA6_7_LC_8_5_3 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_5HZ_RNITRA6_7_LC_8_5_3 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_5HZ_RNITRA6_7_LC_8_5_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_RNITRA6_7_LC_8_5_3  (
            .in0(_gnd_net_),
            .in1(N__2405),
            .in2(_gnd_net_),
            .in3(N__2371),
            .lcout(\LED_Blink_Inst.un1_r_count_5hz_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_1_LC_8_5_5 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_5HZ_1_LC_8_5_5 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_5HZ_1_LC_8_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_1_LC_8_5_5  (
            .in0(N__2393),
            .in1(N__2719),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\LED_Blink_Inst.r_Count_5HZZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4433),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_8_LC_8_5_6 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_5HZ_8_LC_8_5_6 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_5HZ_8_LC_8_5_6 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_8_LC_8_5_6  (
            .in0(N__2515),
            .in1(N__2617),
            .in2(N__2563),
            .in3(N__2378),
            .lcout(\LED_Blink_Inst.r_Count_5HZZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4433),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Toggle_5HZ_LC_8_5_7 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Toggle_5HZ_LC_8_5_7 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Toggle_5HZ_LC_8_5_7 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \LED_Blink_Inst.r_Toggle_5HZ_LC_8_5_7  (
            .in0(N__2618),
            .in1(N__2516),
            .in2(N__2356),
            .in3(N__2556),
            .lcout(o_LED_2_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4433),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_0_LC_8_6_0 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_5HZ_0_LC_8_6_0 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_5HZ_0_LC_8_6_0 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_0_LC_8_6_0  (
            .in0(N__2500),
            .in1(N__2718),
            .in2(N__2612),
            .in3(N__2548),
            .lcout(\LED_Blink_Inst.r_Count_5HZZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4429),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_13_LC_8_6_1 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_5HZ_13_LC_8_6_1 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_5HZ_13_LC_8_6_1 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_13_LC_8_6_1  (
            .in0(N__2595),
            .in1(N__2502),
            .in2(N__2561),
            .in3(N__2339),
            .lcout(\LED_Blink_Inst.r_Count_5HZZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4429),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_RNII1D11_10_LC_8_6_2 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_5HZ_RNII1D11_10_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_5HZ_RNII1D11_10_LC_8_6_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_RNII1D11_10_LC_8_6_2  (
            .in0(N__2333),
            .in1(N__2465),
            .in2(N__2687),
            .in3(N__2320),
            .lcout(),
            .ltout(\LED_Blink_Inst.un1_r_count_5hz_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_RNI5I2E1_3_LC_8_6_3 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_5HZ_RNI5I2E1_3_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_5HZ_RNI5I2E1_3_LC_8_6_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_RNI5I2E1_3_LC_8_6_3  (
            .in0(N__2309),
            .in1(N__2297),
            .in2(N__2285),
            .in3(N__2282),
            .lcout(),
            .ltout(\LED_Blink_Inst.un1_r_count_5hz_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_RNIE3862_11_LC_8_6_4 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_5HZ_RNIE3862_11_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_5HZ_RNIE3862_11_LC_8_6_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_RNIE3862_11_LC_8_6_4  (
            .in0(N__2741),
            .in1(N__2735),
            .in2(N__2723),
            .in3(N__2717),
            .lcout(\LED_Blink_Inst.un1_r_count_5hz_19 ),
            .ltout(\LED_Blink_Inst.un1_r_count_5hz_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_17_LC_8_6_5 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_5HZ_17_LC_8_6_5 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_5HZ_17_LC_8_6_5 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_17_LC_8_6_5  (
            .in0(N__2596),
            .in1(N__2503),
            .in2(N__2696),
            .in3(N__2693),
            .lcout(\LED_Blink_Inst.r_Count_5HZZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4429),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_RNI477S_9_LC_8_6_6 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_5HZ_RNI477S_9_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_5HZ_RNI477S_9_LC_8_6_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_RNI477S_9_LC_8_6_6  (
            .in0(N__2672),
            .in1(N__2660),
            .in2(N__2648),
            .in3(N__2633),
            .lcout(\LED_Blink_Inst.un1_r_count_5hz_15 ),
            .ltout(\LED_Blink_Inst.un1_r_count_5hz_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_5HZ_10_LC_8_6_7 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_5HZ_10_LC_8_6_7 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_5HZ_10_LC_8_6_7 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \LED_Blink_Inst.r_Count_5HZ_10_LC_8_6_7  (
            .in0(N__2544),
            .in1(N__2501),
            .in2(N__2474),
            .in3(N__2471),
            .lcout(\LED_Blink_Inst.r_Count_5HZZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4429),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.un4_r_count_1hz_cry_1_c_LC_8_7_0 .C_ON=1'b1;
    defparam \LED_Blink_Inst.un4_r_count_1hz_cry_1_c_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.un4_r_count_1hz_cry_1_c_LC_8_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \LED_Blink_Inst.un4_r_count_1hz_cry_1_c_LC_8_7_0  (
            .in0(_gnd_net_),
            .in1(N__3171),
            .in2(N__2860),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_7_0_),
            .carryout(\LED_Blink_Inst.un4_r_count_1hz_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_2_LC_8_7_1 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_1HZ_2_LC_8_7_1 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_1HZ_2_LC_8_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_2_LC_8_7_1  (
            .in0(_gnd_net_),
            .in1(N__2821),
            .in2(_gnd_net_),
            .in3(N__2453),
            .lcout(\LED_Blink_Inst.r_Count_1HZZ0Z_2 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_1hz_cry_1 ),
            .carryout(\LED_Blink_Inst.un4_r_count_1hz_cry_2 ),
            .clk(N__4426),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_3_LC_8_7_2 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_1HZ_3_LC_8_7_2 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_1HZ_3_LC_8_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_3_LC_8_7_2  (
            .in0(_gnd_net_),
            .in1(N__2833),
            .in2(_gnd_net_),
            .in3(N__2450),
            .lcout(\LED_Blink_Inst.r_Count_1HZZ0Z_3 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_1hz_cry_2 ),
            .carryout(\LED_Blink_Inst.un4_r_count_1hz_cry_3 ),
            .clk(N__4426),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_4_LC_8_7_3 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_1HZ_4_LC_8_7_3 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_1HZ_4_LC_8_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_4_LC_8_7_3  (
            .in0(_gnd_net_),
            .in1(N__2872),
            .in2(_gnd_net_),
            .in3(N__2447),
            .lcout(\LED_Blink_Inst.r_Count_1HZZ0Z_4 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_1hz_cry_3 ),
            .carryout(\LED_Blink_Inst.un4_r_count_1hz_cry_4 ),
            .clk(N__4426),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_5_LC_8_7_4 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_1HZ_5_LC_8_7_4 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_1HZ_5_LC_8_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_5_LC_8_7_4  (
            .in0(_gnd_net_),
            .in1(N__2911),
            .in2(_gnd_net_),
            .in3(N__2768),
            .lcout(\LED_Blink_Inst.r_Count_1HZZ0Z_5 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_1hz_cry_4 ),
            .carryout(\LED_Blink_Inst.un4_r_count_1hz_cry_5 ),
            .clk(N__4426),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_6_LC_8_7_5 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_1HZ_6_LC_8_7_5 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_1HZ_6_LC_8_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_6_LC_8_7_5  (
            .in0(_gnd_net_),
            .in1(N__2899),
            .in2(_gnd_net_),
            .in3(N__2765),
            .lcout(\LED_Blink_Inst.r_Count_1HZZ0Z_6 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_1hz_cry_5 ),
            .carryout(\LED_Blink_Inst.un4_r_count_1hz_cry_6 ),
            .clk(N__4426),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_7_LC_8_7_6 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_1HZ_7_LC_8_7_6 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_1HZ_7_LC_8_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_7_LC_8_7_6  (
            .in0(_gnd_net_),
            .in1(N__2884),
            .in2(_gnd_net_),
            .in3(N__2762),
            .lcout(\LED_Blink_Inst.r_Count_1HZZ0Z_7 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_1hz_cry_6 ),
            .carryout(\LED_Blink_Inst.un4_r_count_1hz_cry_7 ),
            .clk(N__4426),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_RNO_0_8_LC_8_7_7 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_1HZ_RNO_0_8_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_1HZ_RNO_0_8_LC_8_7_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_RNO_0_8_LC_8_7_7  (
            .in0(_gnd_net_),
            .in1(N__2806),
            .in2(_gnd_net_),
            .in3(N__2759),
            .lcout(\LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_1hz_cry_7 ),
            .carryout(\LED_Blink_Inst.un4_r_count_1hz_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_RNO_0_9_LC_8_8_0 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_1HZ_RNO_0_9_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_1HZ_RNO_0_9_LC_8_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_RNO_0_9_LC_8_8_0  (
            .in0(_gnd_net_),
            .in1(N__3013),
            .in2(_gnd_net_),
            .in3(N__2756),
            .lcout(\LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_8_8_0_),
            .carryout(\LED_Blink_Inst.un4_r_count_1hz_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_10_LC_8_8_1 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_1HZ_10_LC_8_8_1 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_1HZ_10_LC_8_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_10_LC_8_8_1  (
            .in0(_gnd_net_),
            .in1(N__2971),
            .in2(_gnd_net_),
            .in3(N__2753),
            .lcout(\LED_Blink_Inst.r_Count_1HZZ0Z_10 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_1hz_cry_9 ),
            .carryout(\LED_Blink_Inst.un4_r_count_1hz_cry_10 ),
            .clk(N__4422),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_RNO_0_11_LC_8_8_2 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_1HZ_RNO_0_11_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_1HZ_RNO_0_11_LC_8_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_RNO_0_11_LC_8_8_2  (
            .in0(_gnd_net_),
            .in1(N__3148),
            .in2(_gnd_net_),
            .in3(N__2750),
            .lcout(\LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_1hz_cry_10 ),
            .carryout(\LED_Blink_Inst.un4_r_count_1hz_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_RNO_0_12_LC_8_8_3 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_1HZ_RNO_0_12_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_1HZ_RNO_0_12_LC_8_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_RNO_0_12_LC_8_8_3  (
            .in0(_gnd_net_),
            .in1(N__3109),
            .in2(_gnd_net_),
            .in3(N__2747),
            .lcout(\LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_1hz_cry_11 ),
            .carryout(\LED_Blink_Inst.un4_r_count_1hz_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_13_LC_8_8_4 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_1HZ_13_LC_8_8_4 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_1HZ_13_LC_8_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_13_LC_8_8_4  (
            .in0(_gnd_net_),
            .in1(N__2986),
            .in2(_gnd_net_),
            .in3(N__2744),
            .lcout(\LED_Blink_Inst.r_Count_1HZZ0Z_13 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_1hz_cry_12 ),
            .carryout(\LED_Blink_Inst.un4_r_count_1hz_cry_13 ),
            .clk(N__4422),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_14_LC_8_8_5 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_1HZ_14_LC_8_8_5 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_1HZ_14_LC_8_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_14_LC_8_8_5  (
            .in0(_gnd_net_),
            .in1(N__3055),
            .in2(_gnd_net_),
            .in3(N__2795),
            .lcout(\LED_Blink_Inst.r_Count_1HZZ0Z_14 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_1hz_cry_13 ),
            .carryout(\LED_Blink_Inst.un4_r_count_1hz_cry_14 ),
            .clk(N__4422),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_15_LC_8_8_6 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_1HZ_15_LC_8_8_6 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_1HZ_15_LC_8_8_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_15_LC_8_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2956),
            .in3(N__2792),
            .lcout(\LED_Blink_Inst.r_Count_1HZZ0Z_15 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_1hz_cry_14 ),
            .carryout(\LED_Blink_Inst.un4_r_count_1hz_cry_15 ),
            .clk(N__4422),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_RNO_0_16_LC_8_8_7 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_1HZ_RNO_0_16_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_1HZ_RNO_0_16_LC_8_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_RNO_0_16_LC_8_8_7  (
            .in0(_gnd_net_),
            .in1(N__3031),
            .in2(_gnd_net_),
            .in3(N__2789),
            .lcout(\LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_1hz_cry_15 ),
            .carryout(\LED_Blink_Inst.un4_r_count_1hz_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_RNO_0_17_LC_8_9_0 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_1HZ_RNO_0_17_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_1HZ_RNO_0_17_LC_8_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_RNO_0_17_LC_8_9_0  (
            .in0(_gnd_net_),
            .in1(N__3199),
            .in2(_gnd_net_),
            .in3(N__2786),
            .lcout(\LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(bfn_8_9_0_),
            .carryout(\LED_Blink_Inst.un4_r_count_1hz_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_RNO_0_18_LC_8_9_1 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_1HZ_RNO_0_18_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_1HZ_RNO_0_18_LC_8_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_RNO_0_18_LC_8_9_1  (
            .in0(_gnd_net_),
            .in1(N__3226),
            .in2(_gnd_net_),
            .in3(N__2783),
            .lcout(\LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_1hz_cry_17 ),
            .carryout(\LED_Blink_Inst.un4_r_count_1hz_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_19_LC_8_9_2 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_1HZ_19_LC_8_9_2 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_1HZ_19_LC_8_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_19_LC_8_9_2  (
            .in0(_gnd_net_),
            .in1(N__3085),
            .in2(_gnd_net_),
            .in3(N__2780),
            .lcout(\LED_Blink_Inst.r_Count_1HZZ0Z_19 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_1hz_cry_18 ),
            .carryout(\LED_Blink_Inst.un4_r_count_1hz_cry_19 ),
            .clk(N__4427),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_RNO_0_20_LC_8_9_3 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_1HZ_RNO_0_20_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_1HZ_RNO_0_20_LC_8_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_RNO_0_20_LC_8_9_3  (
            .in0(_gnd_net_),
            .in1(N__3239),
            .in2(_gnd_net_),
            .in3(N__2777),
            .lcout(\LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_1hz_cry_19 ),
            .carryout(\LED_Blink_Inst.un4_r_count_1hz_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_RNO_0_21_LC_8_9_4 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_1HZ_RNO_0_21_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_1HZ_RNO_0_21_LC_8_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_RNO_0_21_LC_8_9_4  (
            .in0(_gnd_net_),
            .in1(N__3214),
            .in2(_gnd_net_),
            .in3(N__2774),
            .lcout(\LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_21 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_1hz_cry_20 ),
            .carryout(\LED_Blink_Inst.un4_r_count_1hz_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_22_LC_8_9_5 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_1HZ_22_LC_8_9_5 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_1HZ_22_LC_8_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_22_LC_8_9_5  (
            .in0(_gnd_net_),
            .in1(N__3097),
            .in2(_gnd_net_),
            .in3(N__2771),
            .lcout(\LED_Blink_Inst.r_Count_1HZZ0Z_22 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_1hz_cry_21 ),
            .carryout(\LED_Blink_Inst.un4_r_count_1hz_cry_22 ),
            .clk(N__4427),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_RNO_0_23_LC_8_9_6 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_1HZ_RNO_0_23_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_1HZ_RNO_0_23_LC_8_9_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_RNO_0_23_LC_8_9_6  (
            .in0(_gnd_net_),
            .in1(N__3070),
            .in2(_gnd_net_),
            .in3(N__2996),
            .lcout(),
            .ltout(\LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_23_LC_8_9_7 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_1HZ_23_LC_8_9_7 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_1HZ_23_LC_8_9_7 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_23_LC_8_9_7  (
            .in0(N__3371),
            .in1(N__3283),
            .in2(N__2993),
            .in3(N__3428),
            .lcout(\LED_Blink_Inst.r_Count_1HZZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4427),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_RNI7T7T_10_LC_9_6_3 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_1HZ_RNI7T7T_10_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_1HZ_RNI7T7T_10_LC_9_6_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_RNI7T7T_10_LC_9_6_3  (
            .in0(N__2990),
            .in1(N__2975),
            .in2(N__2960),
            .in3(N__2855),
            .lcout(\LED_Blink_Inst.un1_r_count_1hz_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_8_LC_9_7_0 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_1HZ_8_LC_9_7_0 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_1HZ_8_LC_9_7_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_8_LC_9_7_0  (
            .in0(N__3286),
            .in1(N__3422),
            .in2(N__3373),
            .in3(N__2939),
            .lcout(\LED_Blink_Inst.r_Count_1HZZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4430),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_0_LC_9_7_1 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_1HZ_0_LC_9_7_1 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_1HZ_0_LC_9_7_1 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_0_LC_9_7_1  (
            .in0(N__3420),
            .in1(N__3284),
            .in2(N__3370),
            .in3(N__2856),
            .lcout(\LED_Blink_Inst.r_Count_1HZZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4430),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Toggle_1HZ_LC_9_7_2 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Toggle_1HZ_LC_9_7_2 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Toggle_1HZ_LC_9_7_2 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \LED_Blink_Inst.r_Toggle_1HZ_LC_9_7_2  (
            .in0(N__3287),
            .in1(N__3423),
            .in2(N__2929),
            .in3(N__3346),
            .lcout(o_LED_4_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4430),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_RNI2VI71_4_LC_9_7_3 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_1HZ_RNI2VI71_4_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_1HZ_RNI2VI71_4_LC_9_7_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_RNI2VI71_4_LC_9_7_3  (
            .in0(N__2912),
            .in1(N__2900),
            .in2(N__2888),
            .in3(N__2873),
            .lcout(\LED_Blink_Inst.un1_r_count_1hz_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_1_LC_9_7_4 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_1HZ_1_LC_9_7_4 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_1HZ_1_LC_9_7_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_1_LC_9_7_4  (
            .in0(N__3173),
            .in1(_gnd_net_),
            .in2(N__2861),
            .in3(_gnd_net_),
            .lcout(\LED_Blink_Inst.r_Count_1HZZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4430),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_RNIQMI71_1_LC_9_7_5 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_1HZ_RNIQMI71_1_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_1HZ_RNIQMI71_1_LC_9_7_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_RNIQMI71_1_LC_9_7_5  (
            .in0(N__2834),
            .in1(N__2822),
            .in2(N__2810),
            .in3(N__3172),
            .lcout(\LED_Blink_Inst.un1_r_count_1hz_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_11_LC_9_7_6 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_1HZ_11_LC_9_7_6 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_1HZ_11_LC_9_7_6 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_11_LC_9_7_6  (
            .in0(N__3285),
            .in1(N__3421),
            .in2(N__3158),
            .in3(N__3345),
            .lcout(\LED_Blink_Inst.r_Count_1HZZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4430),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_RNIH78T_11_LC_9_8_0 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_1HZ_RNIH78T_11_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_1HZ_RNIH78T_11_LC_9_8_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_RNIH78T_11_LC_9_8_0  (
            .in0(N__3110),
            .in1(N__3149),
            .in2(N__3035),
            .in3(N__3014),
            .lcout(),
            .ltout(\LED_Blink_Inst.un1_r_count_1hz_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_RNIF0A64_11_LC_9_8_1 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_1HZ_RNIF0A64_11_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_1HZ_RNIF0A64_11_LC_9_8_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_RNIF0A64_11_LC_9_8_1  (
            .in0(N__3188),
            .in1(N__3137),
            .in2(N__3128),
            .in3(N__3125),
            .lcout(\LED_Blink_Inst.un1_r_count_1hz_21 ),
            .ltout(\LED_Blink_Inst.un1_r_count_1hz_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_12_LC_9_8_2 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_1HZ_12_LC_9_8_2 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_1HZ_12_LC_9_8_2 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_12_LC_9_8_2  (
            .in0(N__3350),
            .in1(N__3268),
            .in2(N__3119),
            .in3(N__3116),
            .lcout(\LED_Blink_Inst.r_Count_1HZZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4424),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_RNI45SP_23_LC_9_8_4 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_1HZ_RNI45SP_23_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_1HZ_RNI45SP_23_LC_9_8_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_RNI45SP_23_LC_9_8_4  (
            .in0(N__3098),
            .in1(N__3086),
            .in2(N__3074),
            .in3(N__3056),
            .lcout(\LED_Blink_Inst.un1_r_count_1hz_16 ),
            .ltout(\LED_Blink_Inst.un1_r_count_1hz_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_16_LC_9_8_5 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_1HZ_16_LC_9_8_5 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_1HZ_16_LC_9_8_5 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_16_LC_9_8_5  (
            .in0(N__3369),
            .in1(N__3418),
            .in2(N__3044),
            .in3(N__3041),
            .lcout(\LED_Blink_Inst.r_Count_1HZZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4424),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_9_LC_9_8_6 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_1HZ_9_LC_9_8_6 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_1HZ_9_LC_9_8_6 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_9_LC_9_8_6  (
            .in0(N__3419),
            .in1(N__3269),
            .in2(N__3372),
            .in3(N__3020),
            .lcout(\LED_Blink_Inst.r_Count_1HZZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4424),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_20_LC_9_9_0 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_1HZ_20_LC_9_9_0 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_1HZ_20_LC_9_9_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_20_LC_9_9_0  (
            .in0(N__3281),
            .in1(N__3426),
            .in2(N__3374),
            .in3(N__3002),
            .lcout(\LED_Blink_Inst.r_Count_1HZZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4431),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_18_LC_9_9_3 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_1HZ_18_LC_9_9_3 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_1HZ_18_LC_9_9_3 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_18_LC_9_9_3  (
            .in0(N__3425),
            .in1(N__3280),
            .in2(N__3377),
            .in3(N__3440),
            .lcout(\LED_Blink_Inst.r_Count_1HZZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4431),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_21_LC_9_9_4 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_1HZ_21_LC_9_9_4 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_1HZ_21_LC_9_9_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_21_LC_9_9_4  (
            .in0(N__3282),
            .in1(N__3427),
            .in2(N__3375),
            .in3(N__3434),
            .lcout(\LED_Blink_Inst.r_Count_1HZZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4431),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_17_LC_9_9_5 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_1HZ_17_LC_9_9_5 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_1HZ_17_LC_9_9_5 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_17_LC_9_9_5  (
            .in0(N__3424),
            .in1(N__3383),
            .in2(N__3376),
            .in3(N__3279),
            .lcout(\LED_Blink_Inst.r_Count_1HZZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4431),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_1HZ_RNI23SP_17_LC_9_9_7 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_1HZ_RNI23SP_17_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_1HZ_RNI23SP_17_LC_9_9_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \LED_Blink_Inst.r_Count_1HZ_RNI23SP_17_LC_9_9_7  (
            .in0(N__3238),
            .in1(N__3227),
            .in2(N__3215),
            .in3(N__3200),
            .lcout(\LED_Blink_Inst.un1_r_count_1hz_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.un6_r_count_10hz_cry_1_c_LC_11_3_0 .C_ON=1'b1;
    defparam \LED_Blink_Inst.un6_r_count_10hz_cry_1_c_LC_11_3_0 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.un6_r_count_10hz_cry_1_c_LC_11_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \LED_Blink_Inst.un6_r_count_10hz_cry_1_c_LC_11_3_0  (
            .in0(_gnd_net_),
            .in1(N__4032),
            .in2(N__3680),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_3_0_),
            .carryout(\LED_Blink_Inst.un6_r_count_10hz_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_2_LC_11_3_1 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_10HZ_2_LC_11_3_1 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_10HZ_2_LC_11_3_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_2_LC_11_3_1  (
            .in0(_gnd_net_),
            .in1(N__4045),
            .in2(_gnd_net_),
            .in3(N__3182),
            .lcout(\LED_Blink_Inst.r_Count_10HZZ0Z_2 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un6_r_count_10hz_cry_1 ),
            .carryout(\LED_Blink_Inst.un6_r_count_10hz_cry_2 ),
            .clk(N__4443),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_3_LC_11_3_2 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_10HZ_3_LC_11_3_2 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_10HZ_3_LC_11_3_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_3_LC_11_3_2  (
            .in0(_gnd_net_),
            .in1(N__3691),
            .in2(_gnd_net_),
            .in3(N__3179),
            .lcout(\LED_Blink_Inst.r_Count_10HZZ0Z_3 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un6_r_count_10hz_cry_2 ),
            .carryout(\LED_Blink_Inst.un6_r_count_10hz_cry_3 ),
            .clk(N__4443),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_RNO_0_4_LC_11_3_3 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_10HZ_RNO_0_4_LC_11_3_3 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_10HZ_RNO_0_4_LC_11_3_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_RNO_0_4_LC_11_3_3  (
            .in0(_gnd_net_),
            .in1(N__3658),
            .in2(_gnd_net_),
            .in3(N__3176),
            .lcout(\LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un6_r_count_10hz_cry_3 ),
            .carryout(\LED_Blink_Inst.un6_r_count_10hz_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_5_LC_11_3_4 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_10HZ_5_LC_11_3_4 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_10HZ_5_LC_11_3_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_5_LC_11_3_4  (
            .in0(_gnd_net_),
            .in1(N__3703),
            .in2(_gnd_net_),
            .in3(N__3467),
            .lcout(\LED_Blink_Inst.r_Count_10HZZ0Z_5 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un6_r_count_10hz_cry_4 ),
            .carryout(\LED_Blink_Inst.un6_r_count_10hz_cry_5 ),
            .clk(N__4443),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_RNO_0_6_LC_11_3_5 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_10HZ_RNO_0_6_LC_11_3_5 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_10HZ_RNO_0_6_LC_11_3_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_RNO_0_6_LC_11_3_5  (
            .in0(_gnd_net_),
            .in1(N__3641),
            .in2(_gnd_net_),
            .in3(N__3464),
            .lcout(\LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un6_r_count_10hz_cry_5 ),
            .carryout(\LED_Blink_Inst.un6_r_count_10hz_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_RNO_0_7_LC_11_3_6 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_10HZ_RNO_0_7_LC_11_3_6 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_10HZ_RNO_0_7_LC_11_3_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_RNO_0_7_LC_11_3_6  (
            .in0(_gnd_net_),
            .in1(N__4072),
            .in2(_gnd_net_),
            .in3(N__3461),
            .lcout(\LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un6_r_count_10hz_cry_6 ),
            .carryout(\LED_Blink_Inst.un6_r_count_10hz_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_8_LC_11_3_7 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_10HZ_8_LC_11_3_7 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_10HZ_8_LC_11_3_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_8_LC_11_3_7  (
            .in0(_gnd_net_),
            .in1(N__4006),
            .in2(_gnd_net_),
            .in3(N__3458),
            .lcout(\LED_Blink_Inst.r_Count_10HZZ0Z_8 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un6_r_count_10hz_cry_7 ),
            .carryout(\LED_Blink_Inst.un6_r_count_10hz_cry_8 ),
            .clk(N__4443),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_RNO_0_9_LC_11_4_0 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_10HZ_RNO_0_9_LC_11_4_0 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_10HZ_RNO_0_9_LC_11_4_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_RNO_0_9_LC_11_4_0  (
            .in0(_gnd_net_),
            .in1(N__3961),
            .in2(_gnd_net_),
            .in3(N__3455),
            .lcout(\LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_11_4_0_),
            .carryout(\LED_Blink_Inst.un6_r_count_10hz_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_10_LC_11_4_1 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_10HZ_10_LC_11_4_1 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_10HZ_10_LC_11_4_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_10_LC_11_4_1  (
            .in0(_gnd_net_),
            .in1(N__3994),
            .in2(_gnd_net_),
            .in3(N__3452),
            .lcout(\LED_Blink_Inst.r_Count_10HZZ0Z_10 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un6_r_count_10hz_cry_9 ),
            .carryout(\LED_Blink_Inst.un6_r_count_10hz_cry_10 ),
            .clk(N__4441),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_11_LC_11_4_2 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_10HZ_11_LC_11_4_2 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_10HZ_11_LC_11_4_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_11_LC_11_4_2  (
            .in0(_gnd_net_),
            .in1(N__3577),
            .in2(_gnd_net_),
            .in3(N__3449),
            .lcout(\LED_Blink_Inst.r_Count_10HZZ0Z_11 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un6_r_count_10hz_cry_10 ),
            .carryout(\LED_Blink_Inst.un6_r_count_10hz_cry_11 ),
            .clk(N__4441),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_RNO_0_12_LC_11_4_3 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_10HZ_RNO_0_12_LC_11_4_3 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_10HZ_RNO_0_12_LC_11_4_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_RNO_0_12_LC_11_4_3  (
            .in0(_gnd_net_),
            .in1(N__4084),
            .in2(_gnd_net_),
            .in3(N__3446),
            .lcout(\LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un6_r_count_10hz_cry_11 ),
            .carryout(\LED_Blink_Inst.un6_r_count_10hz_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_13_LC_11_4_4 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_10HZ_13_LC_11_4_4 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_10HZ_13_LC_11_4_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_13_LC_11_4_4  (
            .in0(_gnd_net_),
            .in1(N__3616),
            .in2(_gnd_net_),
            .in3(N__3443),
            .lcout(\LED_Blink_Inst.r_Count_10HZZ0Z_13 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un6_r_count_10hz_cry_12 ),
            .carryout(\LED_Blink_Inst.un6_r_count_10hz_cry_13 ),
            .clk(N__4441),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_14_LC_11_4_5 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_10HZ_14_LC_11_4_5 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_10HZ_14_LC_11_4_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_14_LC_11_4_5  (
            .in0(_gnd_net_),
            .in1(N__3589),
            .in2(_gnd_net_),
            .in3(N__3521),
            .lcout(\LED_Blink_Inst.r_Count_10HZZ0Z_14 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un6_r_count_10hz_cry_13 ),
            .carryout(\LED_Blink_Inst.un6_r_count_10hz_cry_14 ),
            .clk(N__4441),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_15_LC_11_4_6 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_10HZ_15_LC_11_4_6 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_10HZ_15_LC_11_4_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_15_LC_11_4_6  (
            .in0(_gnd_net_),
            .in1(N__3604),
            .in2(_gnd_net_),
            .in3(N__3518),
            .lcout(\LED_Blink_Inst.r_Count_10HZZ0Z_15 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un6_r_count_10hz_cry_14 ),
            .carryout(\LED_Blink_Inst.un6_r_count_10hz_cry_15 ),
            .clk(N__4441),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_RNO_0_16_LC_11_4_7 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_10HZ_RNO_0_16_LC_11_4_7 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_10HZ_RNO_0_16_LC_11_4_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_RNO_0_16_LC_11_4_7  (
            .in0(_gnd_net_),
            .in1(N__4058),
            .in2(_gnd_net_),
            .in3(N__3515),
            .lcout(\LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un6_r_count_10hz_cry_15 ),
            .carryout(\LED_Blink_Inst.un6_r_count_10hz_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_RNO_0_17_LC_11_5_0 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_10HZ_RNO_0_17_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_10HZ_RNO_0_17_LC_11_5_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_RNO_0_17_LC_11_5_0  (
            .in0(_gnd_net_),
            .in1(N__3529),
            .in2(_gnd_net_),
            .in3(N__3512),
            .lcout(\LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(bfn_11_5_0_),
            .carryout(\LED_Blink_Inst.un6_r_count_10hz_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_18_LC_11_5_1 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_10HZ_18_LC_11_5_1 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_10HZ_18_LC_11_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_18_LC_11_5_1  (
            .in0(_gnd_net_),
            .in1(N__3475),
            .in2(_gnd_net_),
            .in3(N__3509),
            .lcout(\LED_Blink_Inst.r_Count_10HZZ0Z_18 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un6_r_count_10hz_cry_17 ),
            .carryout(\LED_Blink_Inst.un6_r_count_10hz_cry_18 ),
            .clk(N__4439),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_19_LC_11_5_2 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_10HZ_19_LC_11_5_2 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_10HZ_19_LC_11_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_19_LC_11_5_2  (
            .in0(_gnd_net_),
            .in1(N__3484),
            .in2(_gnd_net_),
            .in3(N__3506),
            .lcout(\LED_Blink_Inst.r_Count_10HZZ0Z_19 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un6_r_count_10hz_cry_18 ),
            .carryout(\LED_Blink_Inst.un6_r_count_10hz_cry_19 ),
            .clk(N__4439),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_RNO_0_20_LC_11_5_3 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_10HZ_RNO_0_20_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_10HZ_RNO_0_20_LC_11_5_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_RNO_0_20_LC_11_5_3  (
            .in0(_gnd_net_),
            .in1(N__3497),
            .in2(_gnd_net_),
            .in3(N__3503),
            .lcout(),
            .ltout(\LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_20_LC_11_5_4 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_10HZ_20_LC_11_5_4 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_10HZ_20_LC_11_5_4 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_20_LC_11_5_4  (
            .in0(N__3832),
            .in1(N__3945),
            .in2(N__3500),
            .in3(N__3879),
            .lcout(\LED_Blink_Inst.r_Count_10HZZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4439),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_RNI9JA61_20_LC_11_5_5 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_10HZ_RNI9JA61_20_LC_11_5_5 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_10HZ_RNI9JA61_20_LC_11_5_5 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_RNI9JA61_20_LC_11_5_5  (
            .in0(N__3530),
            .in1(N__3496),
            .in2(N__3488),
            .in3(N__3476),
            .lcout(\LED_Blink_Inst.un1_r_count_10hz_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_17_LC_11_5_7 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_10HZ_17_LC_11_5_7 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_10HZ_17_LC_11_5_7 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_17_LC_11_5_7  (
            .in0(N__3878),
            .in1(N__3536),
            .in2(N__3950),
            .in3(N__3833),
            .lcout(\LED_Blink_Inst.r_Count_10HZZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4439),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_1_LC_11_6_0 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_2HZ_1_LC_11_6_0 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_2HZ_1_LC_11_6_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_1_LC_11_6_0  (
            .in0(_gnd_net_),
            .in1(N__3763),
            .in2(_gnd_net_),
            .in3(N__3782),
            .lcout(\LED_Blink_Inst.r_Count_2HZZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4436),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_RNIPIKC_6_LC_11_7_0 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNIPIKC_6_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNIPIKC_6_LC_11_7_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_RNIPIKC_6_LC_11_7_0  (
            .in0(N__4175),
            .in1(N__4190),
            .in2(_gnd_net_),
            .in3(N__3761),
            .lcout(\LED_Blink_Inst.un1_r_count_2hz_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_RNIR7RG_1_LC_11_7_1 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNIR7RG_1_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNIR7RG_1_LC_11_7_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_RNIR7RG_1_LC_11_7_1  (
            .in0(N__3725),
            .in1(N__3781),
            .in2(N__4208),
            .in3(N__3740),
            .lcout(\LED_Blink_Inst.un1_r_count_2hz_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_11_LC_11_7_2 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_2HZ_11_LC_11_7_2 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_2HZ_11_LC_11_7_2 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_11_LC_11_7_2  (
            .in0(N__4578),
            .in1(N__4097),
            .in2(N__4528),
            .in3(N__4643),
            .lcout(\LED_Blink_Inst.r_Count_2HZZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4435),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_0_LC_11_7_3 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_2HZ_0_LC_11_7_3 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_2HZ_0_LC_11_7_3 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_0_LC_11_7_3  (
            .in0(N__3762),
            .in1(N__4641),
            .in2(N__4529),
            .in3(N__4580),
            .lcout(\LED_Blink_Inst.r_Count_2HZZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4435),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_4_LC_11_7_4 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_2HZ_4_LC_11_7_4 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_2HZ_4_LC_11_7_4 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_4_LC_11_7_4  (
            .in0(N__4579),
            .in1(N__4524),
            .in2(N__4220),
            .in3(N__4644),
            .lcout(\LED_Blink_Inst.r_Count_2HZZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4435),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_RNI009U_4_LC_11_7_5 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNI009U_4_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNI009U_4_LC_11_7_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_RNI009U_4_LC_11_7_5  (
            .in0(N__4136),
            .in1(N__4157),
            .in2(N__4112),
            .in3(N__4232),
            .lcout(\LED_Blink_Inst.un1_r_count_2hz_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_9_LC_11_7_6 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_2HZ_9_LC_11_7_6 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_2HZ_9_LC_11_7_6 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_9_LC_11_7_6  (
            .in0(N__4519),
            .in1(N__4645),
            .in2(N__4591),
            .in3(N__4145),
            .lcout(\LED_Blink_Inst.r_Count_2HZZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4435),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_10_LC_11_7_7 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_2HZ_10_LC_11_7_7 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_2HZ_10_LC_11_7_7 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_10_LC_11_7_7  (
            .in0(N__4642),
            .in1(N__4520),
            .in2(N__4124),
            .in3(N__4584),
            .lcout(\LED_Blink_Inst.r_Count_2HZZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4435),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_16_LC_11_8_0 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_2HZ_16_LC_11_8_0 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_2HZ_16_LC_11_8_0 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_16_LC_11_8_0  (
            .in0(N__4638),
            .in1(N__4573),
            .in2(N__4298),
            .in3(N__4513),
            .lcout(\LED_Blink_Inst.r_Count_2HZZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4432),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_20_LC_11_8_1 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_2HZ_20_LC_11_8_1 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_2HZ_20_LC_11_8_1 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_20_LC_11_8_1  (
            .in0(N__4511),
            .in1(N__4640),
            .in2(N__4590),
            .in3(N__4241),
            .lcout(\LED_Blink_Inst.r_Count_2HZZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4432),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_19_LC_11_8_2 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_2HZ_19_LC_11_8_2 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_2HZ_19_LC_11_8_2 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_19_LC_11_8_2  (
            .in0(N__4639),
            .in1(N__4574),
            .in2(N__4265),
            .in3(N__4514),
            .lcout(\LED_Blink_Inst.r_Count_2HZZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4432),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_RNI7QMB1_12_LC_11_8_3 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNI7QMB1_12_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNI7QMB1_12_LC_11_8_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_RNI7QMB1_12_LC_11_8_3  (
            .in0(N__4310),
            .in1(N__4334),
            .in2(N__4682),
            .in3(N__4367),
            .lcout(),
            .ltout(\LED_Blink_Inst.un1_r_count_2hz_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_RNIRKF73_1_LC_11_8_4 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNIRKF73_1_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNIRKF73_1_LC_11_8_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_RNIRKF73_1_LC_11_8_4  (
            .in0(N__3566),
            .in1(N__3560),
            .in2(N__3554),
            .in3(N__3551),
            .lcout(\LED_Blink_Inst.un1_r_count_2hz_20 ),
            .ltout(\LED_Blink_Inst.un1_r_count_2hz_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_14_LC_11_8_5 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_2HZ_14_LC_11_8_5 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_2HZ_14_LC_11_8_5 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_14_LC_11_8_5  (
            .in0(N__4571),
            .in1(N__4637),
            .in2(N__3545),
            .in3(N__4322),
            .lcout(\LED_Blink_Inst.r_Count_2HZZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4432),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_12_LC_11_8_6 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_2HZ_12_LC_11_8_6 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_2HZ_12_LC_11_8_6 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_12_LC_11_8_6  (
            .in0(N__4636),
            .in1(N__4572),
            .in2(N__4355),
            .in3(N__4512),
            .lcout(\LED_Blink_Inst.r_Count_2HZZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4432),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_RNI9UOB1_22_LC_11_8_7 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNI9UOB1_22_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNI9UOB1_22_LC_11_8_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_RNI9UOB1_22_LC_11_8_7  (
            .in0(N__4661),
            .in1(N__4253),
            .in2(N__4757),
            .in3(N__4277),
            .lcout(\LED_Blink_Inst.un1_r_count_2hz_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_0_LC_12_3_0 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_10HZ_0_LC_12_3_0 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_10HZ_0_LC_12_3_0 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_0_LC_12_3_0  (
            .in0(N__3678),
            .in1(N__3885),
            .in2(N__3948),
            .in3(N__3830),
            .lcout(\LED_Blink_Inst.r_Count_10HZZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4445),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_7_LC_12_3_1 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_10HZ_7_LC_12_3_1 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_10HZ_7_LC_12_3_1 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_7_LC_12_3_1  (
            .in0(N__3829),
            .in1(N__3940),
            .in2(N__3893),
            .in3(N__3542),
            .lcout(\LED_Blink_Inst.r_Count_10HZZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4445),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_4_LC_12_3_2 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_10HZ_4_LC_12_3_2 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_10HZ_4_LC_12_3_2 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_4_LC_12_3_2  (
            .in0(N__3884),
            .in1(N__3710),
            .in2(N__3949),
            .in3(N__3831),
            .lcout(\LED_Blink_Inst.r_Count_10HZZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4445),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_RNI1U1B_3_LC_12_3_3 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_10HZ_RNI1U1B_3_LC_12_3_3 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_10HZ_RNI1U1B_3_LC_12_3_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_RNI1U1B_3_LC_12_3_3  (
            .in0(N__3704),
            .in1(N__3692),
            .in2(_gnd_net_),
            .in3(N__3677),
            .lcout(\LED_Blink_Inst.un1_r_count_10hz_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_1_LC_12_3_4 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_10HZ_1_LC_12_3_4 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_10HZ_1_LC_12_3_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_1_LC_12_3_4  (
            .in0(N__3679),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4034),
            .lcout(\LED_Blink_Inst.r_Count_10HZZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4445),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_RNIG3C7_4_LC_12_3_5 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_10HZ_RNIG3C7_4_LC_12_3_5 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_10HZ_RNIG3C7_4_LC_12_3_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_RNIG3C7_4_LC_12_3_5  (
            .in0(_gnd_net_),
            .in1(N__3659),
            .in2(_gnd_net_),
            .in3(N__3640),
            .lcout(\LED_Blink_Inst.un1_r_count_10hz_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_6_LC_12_3_7 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_10HZ_6_LC_12_3_7 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_10HZ_6_LC_12_3_7 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_6_LC_12_3_7  (
            .in0(N__3828),
            .in1(N__3939),
            .in2(N__3892),
            .in3(N__3647),
            .lcout(\LED_Blink_Inst.r_Count_10HZZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4445),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_16_LC_12_4_0 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_10HZ_16_LC_12_4_0 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_10HZ_16_LC_12_4_0 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_16_LC_12_4_0  (
            .in0(N__3881),
            .in1(N__3629),
            .in2(N__3947),
            .in3(N__3835),
            .lcout(\LED_Blink_Inst.r_Count_10HZZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4444),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_12_LC_12_4_2 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_10HZ_12_LC_12_4_2 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_10HZ_12_LC_12_4_2 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_12_LC_12_4_2  (
            .in0(N__3880),
            .in1(N__3623),
            .in2(N__3946),
            .in3(N__3834),
            .lcout(\LED_Blink_Inst.r_Count_10HZZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4444),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_RNIT5961_11_LC_12_4_3 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_10HZ_RNIT5961_11_LC_12_4_3 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_10HZ_RNIT5961_11_LC_12_4_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_RNIT5961_11_LC_12_4_3  (
            .in0(N__3617),
            .in1(N__3605),
            .in2(N__3593),
            .in3(N__3578),
            .lcout(\LED_Blink_Inst.un1_r_count_10hz_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_RNI6UGQ_7_LC_12_4_4 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_10HZ_RNI6UGQ_7_LC_12_4_4 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_10HZ_RNI6UGQ_7_LC_12_4_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_RNI6UGQ_7_LC_12_4_4  (
            .in0(N__4085),
            .in1(N__3962),
            .in2(N__4073),
            .in3(N__4057),
            .lcout(),
            .ltout(\LED_Blink_Inst.un1_r_count_10hz_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_RNIVT891_1_LC_12_4_5 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_10HZ_RNIVT891_1_LC_12_4_5 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_10HZ_RNIVT891_1_LC_12_4_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_RNIVT891_1_LC_12_4_5  (
            .in0(N__4046),
            .in1(N__4033),
            .in2(N__4016),
            .in3(N__4013),
            .lcout(),
            .ltout(\LED_Blink_Inst.un1_r_count_10hz_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_RNIV6J12_8_LC_12_4_6 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_10HZ_RNIV6J12_8_LC_12_4_6 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_10HZ_RNIV6J12_8_LC_12_4_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_RNIV6J12_8_LC_12_4_6  (
            .in0(N__4007),
            .in1(N__3995),
            .in2(N__3983),
            .in3(N__3980),
            .lcout(\LED_Blink_Inst.un1_r_count_10hz_18 ),
            .ltout(\LED_Blink_Inst.un1_r_count_10hz_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_10HZ_9_LC_12_4_7 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_10HZ_9_LC_12_4_7 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_10HZ_9_LC_12_4_7 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \LED_Blink_Inst.r_Count_10HZ_9_LC_12_4_7  (
            .in0(N__3883),
            .in1(N__3971),
            .in2(N__3965),
            .in3(N__3932),
            .lcout(\LED_Blink_Inst.r_Count_10HZZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4444),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Toggle_10HZ_LC_12_5_4 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Toggle_10HZ_LC_12_5_4 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Toggle_10HZ_LC_12_5_4 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \LED_Blink_Inst.r_Toggle_10HZ_LC_12_5_4  (
            .in0(N__3941),
            .in1(N__3882),
            .in2(N__3797),
            .in3(N__3836),
            .lcout(o_LED_1_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4442),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.un4_r_count_2hz_cry_1_c_LC_12_6_0 .C_ON=1'b1;
    defparam \LED_Blink_Inst.un4_r_count_2hz_cry_1_c_LC_12_6_0 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.un4_r_count_2hz_cry_1_c_LC_12_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \LED_Blink_Inst.un4_r_count_2hz_cry_1_c_LC_12_6_0  (
            .in0(_gnd_net_),
            .in1(N__3780),
            .in2(N__3764),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_6_0_),
            .carryout(\LED_Blink_Inst.un4_r_count_2hz_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_2_LC_12_6_1 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_2HZ_2_LC_12_6_1 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_2HZ_2_LC_12_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_2_LC_12_6_1  (
            .in0(_gnd_net_),
            .in1(N__3739),
            .in2(_gnd_net_),
            .in3(N__3728),
            .lcout(\LED_Blink_Inst.r_Count_2HZZ0Z_2 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_2hz_cry_1 ),
            .carryout(\LED_Blink_Inst.un4_r_count_2hz_cry_2 ),
            .clk(N__4440),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_3_LC_12_6_2 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_2HZ_3_LC_12_6_2 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_2HZ_3_LC_12_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_3_LC_12_6_2  (
            .in0(_gnd_net_),
            .in1(N__3724),
            .in2(_gnd_net_),
            .in3(N__3713),
            .lcout(\LED_Blink_Inst.r_Count_2HZZ0Z_3 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_2hz_cry_2 ),
            .carryout(\LED_Blink_Inst.un4_r_count_2hz_cry_3 ),
            .clk(N__4440),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_4_LC_12_6_3 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_4_LC_12_6_3 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_4_LC_12_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_RNO_0_4_LC_12_6_3  (
            .in0(_gnd_net_),
            .in1(N__4231),
            .in2(_gnd_net_),
            .in3(N__4211),
            .lcout(\LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_2hz_cry_3 ),
            .carryout(\LED_Blink_Inst.un4_r_count_2hz_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_5_LC_12_6_4 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_2HZ_5_LC_12_6_4 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_2HZ_5_LC_12_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_5_LC_12_6_4  (
            .in0(_gnd_net_),
            .in1(N__4204),
            .in2(_gnd_net_),
            .in3(N__4193),
            .lcout(\LED_Blink_Inst.r_Count_2HZZ0Z_5 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_2hz_cry_4 ),
            .carryout(\LED_Blink_Inst.un4_r_count_2hz_cry_5 ),
            .clk(N__4440),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_6_LC_12_6_5 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_2HZ_6_LC_12_6_5 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_2HZ_6_LC_12_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_6_LC_12_6_5  (
            .in0(_gnd_net_),
            .in1(N__4189),
            .in2(_gnd_net_),
            .in3(N__4178),
            .lcout(\LED_Blink_Inst.r_Count_2HZZ0Z_6 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_2hz_cry_5 ),
            .carryout(\LED_Blink_Inst.un4_r_count_2hz_cry_6 ),
            .clk(N__4440),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_7_LC_12_6_6 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_2HZ_7_LC_12_6_6 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_2HZ_7_LC_12_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_7_LC_12_6_6  (
            .in0(_gnd_net_),
            .in1(N__4174),
            .in2(_gnd_net_),
            .in3(N__4163),
            .lcout(\LED_Blink_Inst.r_Count_2HZZ0Z_7 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_2hz_cry_6 ),
            .carryout(\LED_Blink_Inst.un4_r_count_2hz_cry_7 ),
            .clk(N__4440),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_8_LC_12_6_7 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_2HZ_8_LC_12_6_7 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_2HZ_8_LC_12_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_8_LC_12_6_7  (
            .in0(_gnd_net_),
            .in1(N__4702),
            .in2(_gnd_net_),
            .in3(N__4160),
            .lcout(\LED_Blink_Inst.r_Count_2HZZ0Z_8 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_2hz_cry_7 ),
            .carryout(\LED_Blink_Inst.un4_r_count_2hz_cry_8 ),
            .clk(N__4440),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_9_LC_12_7_0 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_9_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_9_LC_12_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_RNO_0_9_LC_12_7_0  (
            .in0(_gnd_net_),
            .in1(N__4156),
            .in2(_gnd_net_),
            .in3(N__4139),
            .lcout(\LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_12_7_0_),
            .carryout(\LED_Blink_Inst.un4_r_count_2hz_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_10_LC_12_7_1 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_10_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_10_LC_12_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_RNO_0_10_LC_12_7_1  (
            .in0(_gnd_net_),
            .in1(N__4135),
            .in2(_gnd_net_),
            .in3(N__4115),
            .lcout(\LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_2hz_cry_9 ),
            .carryout(\LED_Blink_Inst.un4_r_count_2hz_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_11_LC_12_7_2 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_11_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_11_LC_12_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_RNO_0_11_LC_12_7_2  (
            .in0(_gnd_net_),
            .in1(N__4108),
            .in2(_gnd_net_),
            .in3(N__4088),
            .lcout(\LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_2hz_cry_10 ),
            .carryout(\LED_Blink_Inst.un4_r_count_2hz_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_12_LC_12_7_3 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_12_LC_12_7_3 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_12_LC_12_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_RNO_0_12_LC_12_7_3  (
            .in0(_gnd_net_),
            .in1(N__4366),
            .in2(_gnd_net_),
            .in3(N__4340),
            .lcout(\LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_2hz_cry_11 ),
            .carryout(\LED_Blink_Inst.un4_r_count_2hz_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_13_LC_12_7_4 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_2HZ_13_LC_12_7_4 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_2HZ_13_LC_12_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_13_LC_12_7_4  (
            .in0(_gnd_net_),
            .in1(N__4729),
            .in2(_gnd_net_),
            .in3(N__4337),
            .lcout(\LED_Blink_Inst.r_Count_2HZZ0Z_13 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_2hz_cry_12 ),
            .carryout(\LED_Blink_Inst.un4_r_count_2hz_cry_13 ),
            .clk(N__4437),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_14_LC_12_7_5 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_14_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_14_LC_12_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_RNO_0_14_LC_12_7_5  (
            .in0(_gnd_net_),
            .in1(N__4333),
            .in2(_gnd_net_),
            .in3(N__4316),
            .lcout(\LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_2hz_cry_13 ),
            .carryout(\LED_Blink_Inst.un4_r_count_2hz_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_15_LC_12_7_6 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_2HZ_15_LC_12_7_6 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_2HZ_15_LC_12_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_15_LC_12_7_6  (
            .in0(_gnd_net_),
            .in1(N__4741),
            .in2(_gnd_net_),
            .in3(N__4313),
            .lcout(\LED_Blink_Inst.r_Count_2HZZ0Z_15 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_2hz_cry_14 ),
            .carryout(\LED_Blink_Inst.un4_r_count_2hz_cry_15 ),
            .clk(N__4437),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_16_LC_12_7_7 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_16_LC_12_7_7 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_16_LC_12_7_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_RNO_0_16_LC_12_7_7  (
            .in0(_gnd_net_),
            .in1(N__4309),
            .in2(_gnd_net_),
            .in3(N__4286),
            .lcout(\LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_2hz_cry_15 ),
            .carryout(\LED_Blink_Inst.un4_r_count_2hz_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_17_LC_12_8_0 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_17_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_17_LC_12_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_RNO_0_17_LC_12_8_0  (
            .in0(_gnd_net_),
            .in1(N__4678),
            .in2(_gnd_net_),
            .in3(N__4283),
            .lcout(\LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(bfn_12_8_0_),
            .carryout(\LED_Blink_Inst.un4_r_count_2hz_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_18_LC_12_8_1 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_18_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_18_LC_12_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_RNO_0_18_LC_12_8_1  (
            .in0(_gnd_net_),
            .in1(N__4660),
            .in2(_gnd_net_),
            .in3(N__4280),
            .lcout(\LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_2hz_cry_17 ),
            .carryout(\LED_Blink_Inst.un4_r_count_2hz_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_19_LC_12_8_2 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_19_LC_12_8_2 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_19_LC_12_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_RNO_0_19_LC_12_8_2  (
            .in0(_gnd_net_),
            .in1(N__4276),
            .in2(_gnd_net_),
            .in3(N__4256),
            .lcout(\LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_2hz_cry_18 ),
            .carryout(\LED_Blink_Inst.un4_r_count_2hz_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_20_LC_12_8_3 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_20_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_20_LC_12_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_RNO_0_20_LC_12_8_3  (
            .in0(_gnd_net_),
            .in1(N__4252),
            .in2(_gnd_net_),
            .in3(N__4235),
            .lcout(\LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_2hz_cry_19 ),
            .carryout(\LED_Blink_Inst.un4_r_count_2hz_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_21_LC_12_8_4 .C_ON=1'b1;
    defparam \LED_Blink_Inst.r_Count_2HZ_21_LC_12_8_4 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_2HZ_21_LC_12_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_21_LC_12_8_4  (
            .in0(_gnd_net_),
            .in1(N__4714),
            .in2(_gnd_net_),
            .in3(N__4766),
            .lcout(\LED_Blink_Inst.r_Count_2HZZ0Z_21 ),
            .ltout(),
            .carryin(\LED_Blink_Inst.un4_r_count_2hz_cry_20 ),
            .carryout(\LED_Blink_Inst.un4_r_count_2hz_cry_21 ),
            .clk(N__4434),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_22_LC_12_8_5 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_22_LC_12_8_5 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNO_0_22_LC_12_8_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_RNO_0_22_LC_12_8_5  (
            .in0(_gnd_net_),
            .in1(N__4756),
            .in2(_gnd_net_),
            .in3(N__4763),
            .lcout(),
            .ltout(\LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_22_LC_12_8_6 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_2HZ_22_LC_12_8_6 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_2HZ_22_LC_12_8_6 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_22_LC_12_8_6  (
            .in0(N__4570),
            .in1(N__4646),
            .in2(N__4760),
            .in3(N__4518),
            .lcout(\LED_Blink_Inst.r_Count_2HZZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4434),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_RNILV051_8_LC_12_8_7 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNILV051_8_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \LED_Blink_Inst.r_Count_2HZ_RNILV051_8_LC_12_8_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_RNILV051_8_LC_12_8_7  (
            .in0(N__4742),
            .in1(N__4730),
            .in2(N__4718),
            .in3(N__4706),
            .lcout(\LED_Blink_Inst.un1_r_count_2hz_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_17_LC_12_9_0 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_2HZ_17_LC_12_9_0 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_2HZ_17_LC_12_9_0 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_17_LC_12_9_0  (
            .in0(N__4647),
            .in1(N__4586),
            .in2(N__4691),
            .in3(N__4516),
            .lcout(\LED_Blink_Inst.r_Count_2HZZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4438),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Count_2HZ_18_LC_12_9_3 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Count_2HZ_18_LC_12_9_3 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Count_2HZ_18_LC_12_9_3 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \LED_Blink_Inst.r_Count_2HZ_18_LC_12_9_3  (
            .in0(N__4515),
            .in1(N__4648),
            .in2(N__4592),
            .in3(N__4667),
            .lcout(\LED_Blink_Inst.r_Count_2HZZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4438),
            .ce(),
            .sr(_gnd_net_));
    defparam \LED_Blink_Inst.r_Toggle_2HZ_LC_12_9_6 .C_ON=1'b0;
    defparam \LED_Blink_Inst.r_Toggle_2HZ_LC_12_9_6 .SEQ_MODE=4'b1000;
    defparam \LED_Blink_Inst.r_Toggle_2HZ_LC_12_9_6 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \LED_Blink_Inst.r_Toggle_2HZ_LC_12_9_6  (
            .in0(N__4649),
            .in1(N__4585),
            .in2(N__4462),
            .in3(N__4517),
            .lcout(o_LED_3_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4438),
            .ce(),
            .sr(_gnd_net_));
endmodule // LED_Blink_Top_Module
