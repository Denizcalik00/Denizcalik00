-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Feb 19 2025 16:49:25

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "LED_Blink_Top_Module" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of LED_Blink_Top_Module
entity LED_Blink_Top_Module is
port (
    o_LED_3 : out std_logic;
    o_LED_1 : out std_logic;
    i_Clk : in std_logic;
    o_LED_4 : out std_logic;
    o_LED_2 : out std_logic);
end LED_Blink_Top_Module;

-- Architecture of LED_Blink_Top_Module
-- View name is \INTERFACE\
architecture \INTERFACE\ of LED_Blink_Top_Module is

signal \N__4823\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4801\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4784\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4756\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4730\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4691\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4675\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4644\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4641\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4603\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4590\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4579\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4573\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4570\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4552\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4528\ : std_logic;
signal \N__4525\ : std_logic;
signal \N__4524\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4519\ : std_logic;
signal \N__4518\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4515\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4512\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4506\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4459\ : std_logic;
signal \N__4456\ : std_logic;
signal \N__4453\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4445\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4437\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4433\ : std_logic;
signal \N__4432\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4423\ : std_logic;
signal \N__4422\ : std_logic;
signal \N__4373\ : std_logic;
signal \N__4370\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4366\ : std_logic;
signal \N__4363\ : std_logic;
signal \N__4360\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4346\ : std_logic;
signal \N__4343\ : std_logic;
signal \N__4340\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4334\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4322\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4306\ : std_logic;
signal \N__4303\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4289\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4283\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4277\ : std_logic;
signal \N__4276\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4270\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4252\ : std_logic;
signal \N__4249\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4235\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4231\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4225\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4211\ : std_logic;
signal \N__4208\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4201\ : std_logic;
signal \N__4198\ : std_logic;
signal \N__4193\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4189\ : std_logic;
signal \N__4186\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4178\ : std_logic;
signal \N__4175\ : std_logic;
signal \N__4174\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4168\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4156\ : std_logic;
signal \N__4153\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4145\ : std_logic;
signal \N__4142\ : std_logic;
signal \N__4139\ : std_logic;
signal \N__4136\ : std_logic;
signal \N__4135\ : std_logic;
signal \N__4132\ : std_logic;
signal \N__4129\ : std_logic;
signal \N__4124\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4108\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4084\ : std_logic;
signal \N__4081\ : std_logic;
signal \N__4078\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4072\ : std_logic;
signal \N__4069\ : std_logic;
signal \N__4066\ : std_logic;
signal \N__4063\ : std_logic;
signal \N__4058\ : std_logic;
signal \N__4057\ : std_logic;
signal \N__4054\ : std_logic;
signal \N__4051\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4045\ : std_logic;
signal \N__4042\ : std_logic;
signal \N__4039\ : std_logic;
signal \N__4034\ : std_logic;
signal \N__4033\ : std_logic;
signal \N__4032\ : std_logic;
signal \N__4029\ : std_logic;
signal \N__4026\ : std_logic;
signal \N__4023\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4013\ : std_logic;
signal \N__4010\ : std_logic;
signal \N__4007\ : std_logic;
signal \N__4006\ : std_logic;
signal \N__4003\ : std_logic;
signal \N__4000\ : std_logic;
signal \N__3995\ : std_logic;
signal \N__3994\ : std_logic;
signal \N__3991\ : std_logic;
signal \N__3988\ : std_logic;
signal \N__3983\ : std_logic;
signal \N__3980\ : std_logic;
signal \N__3977\ : std_logic;
signal \N__3974\ : std_logic;
signal \N__3971\ : std_logic;
signal \N__3968\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3962\ : std_logic;
signal \N__3961\ : std_logic;
signal \N__3958\ : std_logic;
signal \N__3955\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3949\ : std_logic;
signal \N__3948\ : std_logic;
signal \N__3947\ : std_logic;
signal \N__3946\ : std_logic;
signal \N__3945\ : std_logic;
signal \N__3942\ : std_logic;
signal \N__3941\ : std_logic;
signal \N__3940\ : std_logic;
signal \N__3939\ : std_logic;
signal \N__3936\ : std_logic;
signal \N__3933\ : std_logic;
signal \N__3932\ : std_logic;
signal \N__3929\ : std_logic;
signal \N__3926\ : std_logic;
signal \N__3921\ : std_logic;
signal \N__3918\ : std_logic;
signal \N__3909\ : std_logic;
signal \N__3902\ : std_logic;
signal \N__3893\ : std_logic;
signal \N__3892\ : std_logic;
signal \N__3889\ : std_logic;
signal \N__3886\ : std_logic;
signal \N__3885\ : std_logic;
signal \N__3884\ : std_logic;
signal \N__3883\ : std_logic;
signal \N__3882\ : std_logic;
signal \N__3881\ : std_logic;
signal \N__3880\ : std_logic;
signal \N__3879\ : std_logic;
signal \N__3878\ : std_logic;
signal \N__3871\ : std_logic;
signal \N__3868\ : std_logic;
signal \N__3865\ : std_logic;
signal \N__3862\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3852\ : std_logic;
signal \N__3847\ : std_logic;
signal \N__3836\ : std_logic;
signal \N__3835\ : std_logic;
signal \N__3834\ : std_logic;
signal \N__3833\ : std_logic;
signal \N__3832\ : std_logic;
signal \N__3831\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3829\ : std_logic;
signal \N__3828\ : std_logic;
signal \N__3825\ : std_logic;
signal \N__3820\ : std_logic;
signal \N__3815\ : std_logic;
signal \N__3806\ : std_logic;
signal \N__3797\ : std_logic;
signal \N__3796\ : std_logic;
signal \N__3793\ : std_logic;
signal \N__3790\ : std_logic;
signal \N__3787\ : std_logic;
signal \N__3782\ : std_logic;
signal \N__3781\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3774\ : std_logic;
signal \N__3771\ : std_logic;
signal \N__3764\ : std_logic;
signal \N__3763\ : std_logic;
signal \N__3762\ : std_logic;
signal \N__3761\ : std_logic;
signal \N__3758\ : std_logic;
signal \N__3755\ : std_logic;
signal \N__3750\ : std_logic;
signal \N__3747\ : std_logic;
signal \N__3740\ : std_logic;
signal \N__3739\ : std_logic;
signal \N__3736\ : std_logic;
signal \N__3733\ : std_logic;
signal \N__3728\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3724\ : std_logic;
signal \N__3721\ : std_logic;
signal \N__3718\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3710\ : std_logic;
signal \N__3707\ : std_logic;
signal \N__3704\ : std_logic;
signal \N__3703\ : std_logic;
signal \N__3700\ : std_logic;
signal \N__3697\ : std_logic;
signal \N__3692\ : std_logic;
signal \N__3691\ : std_logic;
signal \N__3688\ : std_logic;
signal \N__3685\ : std_logic;
signal \N__3680\ : std_logic;
signal \N__3679\ : std_logic;
signal \N__3678\ : std_logic;
signal \N__3677\ : std_logic;
signal \N__3674\ : std_logic;
signal \N__3667\ : std_logic;
signal \N__3664\ : std_logic;
signal \N__3659\ : std_logic;
signal \N__3658\ : std_logic;
signal \N__3655\ : std_logic;
signal \N__3652\ : std_logic;
signal \N__3647\ : std_logic;
signal \N__3644\ : std_logic;
signal \N__3641\ : std_logic;
signal \N__3640\ : std_logic;
signal \N__3637\ : std_logic;
signal \N__3634\ : std_logic;
signal \N__3629\ : std_logic;
signal \N__3626\ : std_logic;
signal \N__3623\ : std_logic;
signal \N__3620\ : std_logic;
signal \N__3617\ : std_logic;
signal \N__3616\ : std_logic;
signal \N__3613\ : std_logic;
signal \N__3610\ : std_logic;
signal \N__3605\ : std_logic;
signal \N__3604\ : std_logic;
signal \N__3601\ : std_logic;
signal \N__3598\ : std_logic;
signal \N__3593\ : std_logic;
signal \N__3590\ : std_logic;
signal \N__3589\ : std_logic;
signal \N__3586\ : std_logic;
signal \N__3583\ : std_logic;
signal \N__3578\ : std_logic;
signal \N__3577\ : std_logic;
signal \N__3574\ : std_logic;
signal \N__3571\ : std_logic;
signal \N__3566\ : std_logic;
signal \N__3563\ : std_logic;
signal \N__3560\ : std_logic;
signal \N__3557\ : std_logic;
signal \N__3554\ : std_logic;
signal \N__3551\ : std_logic;
signal \N__3548\ : std_logic;
signal \N__3545\ : std_logic;
signal \N__3542\ : std_logic;
signal \N__3539\ : std_logic;
signal \N__3536\ : std_logic;
signal \N__3533\ : std_logic;
signal \N__3530\ : std_logic;
signal \N__3529\ : std_logic;
signal \N__3524\ : std_logic;
signal \N__3521\ : std_logic;
signal \N__3518\ : std_logic;
signal \N__3515\ : std_logic;
signal \N__3512\ : std_logic;
signal \N__3509\ : std_logic;
signal \N__3506\ : std_logic;
signal \N__3503\ : std_logic;
signal \N__3500\ : std_logic;
signal \N__3497\ : std_logic;
signal \N__3496\ : std_logic;
signal \N__3491\ : std_logic;
signal \N__3488\ : std_logic;
signal \N__3485\ : std_logic;
signal \N__3484\ : std_logic;
signal \N__3479\ : std_logic;
signal \N__3476\ : std_logic;
signal \N__3475\ : std_logic;
signal \N__3470\ : std_logic;
signal \N__3467\ : std_logic;
signal \N__3464\ : std_logic;
signal \N__3461\ : std_logic;
signal \N__3458\ : std_logic;
signal \N__3455\ : std_logic;
signal \N__3452\ : std_logic;
signal \N__3449\ : std_logic;
signal \N__3446\ : std_logic;
signal \N__3443\ : std_logic;
signal \N__3440\ : std_logic;
signal \N__3437\ : std_logic;
signal \N__3434\ : std_logic;
signal \N__3431\ : std_logic;
signal \N__3428\ : std_logic;
signal \N__3427\ : std_logic;
signal \N__3426\ : std_logic;
signal \N__3425\ : std_logic;
signal \N__3424\ : std_logic;
signal \N__3423\ : std_logic;
signal \N__3422\ : std_logic;
signal \N__3421\ : std_logic;
signal \N__3420\ : std_logic;
signal \N__3419\ : std_logic;
signal \N__3418\ : std_logic;
signal \N__3415\ : std_logic;
signal \N__3406\ : std_logic;
signal \N__3397\ : std_logic;
signal \N__3392\ : std_logic;
signal \N__3383\ : std_logic;
signal \N__3380\ : std_logic;
signal \N__3377\ : std_logic;
signal \N__3376\ : std_logic;
signal \N__3375\ : std_logic;
signal \N__3374\ : std_logic;
signal \N__3373\ : std_logic;
signal \N__3372\ : std_logic;
signal \N__3371\ : std_logic;
signal \N__3370\ : std_logic;
signal \N__3369\ : std_logic;
signal \N__3366\ : std_logic;
signal \N__3363\ : std_logic;
signal \N__3360\ : std_logic;
signal \N__3357\ : std_logic;
signal \N__3354\ : std_logic;
signal \N__3351\ : std_logic;
signal \N__3350\ : std_logic;
signal \N__3347\ : std_logic;
signal \N__3346\ : std_logic;
signal \N__3345\ : std_logic;
signal \N__3342\ : std_logic;
signal \N__3339\ : std_logic;
signal \N__3334\ : std_logic;
signal \N__3329\ : std_logic;
signal \N__3326\ : std_logic;
signal \N__3321\ : std_logic;
signal \N__3318\ : std_logic;
signal \N__3311\ : std_logic;
signal \N__3308\ : std_logic;
signal \N__3303\ : std_logic;
signal \N__3296\ : std_logic;
signal \N__3287\ : std_logic;
signal \N__3286\ : std_logic;
signal \N__3285\ : std_logic;
signal \N__3284\ : std_logic;
signal \N__3283\ : std_logic;
signal \N__3282\ : std_logic;
signal \N__3281\ : std_logic;
signal \N__3280\ : std_logic;
signal \N__3279\ : std_logic;
signal \N__3270\ : std_logic;
signal \N__3269\ : std_logic;
signal \N__3268\ : std_logic;
signal \N__3265\ : std_logic;
signal \N__3256\ : std_logic;
signal \N__3253\ : std_logic;
signal \N__3248\ : std_logic;
signal \N__3239\ : std_logic;
signal \N__3238\ : std_logic;
signal \N__3235\ : std_logic;
signal \N__3232\ : std_logic;
signal \N__3227\ : std_logic;
signal \N__3226\ : std_logic;
signal \N__3223\ : std_logic;
signal \N__3220\ : std_logic;
signal \N__3215\ : std_logic;
signal \N__3214\ : std_logic;
signal \N__3211\ : std_logic;
signal \N__3208\ : std_logic;
signal \N__3205\ : std_logic;
signal \N__3200\ : std_logic;
signal \N__3199\ : std_logic;
signal \N__3196\ : std_logic;
signal \N__3193\ : std_logic;
signal \N__3188\ : std_logic;
signal \N__3185\ : std_logic;
signal \N__3182\ : std_logic;
signal \N__3179\ : std_logic;
signal \N__3176\ : std_logic;
signal \N__3173\ : std_logic;
signal \N__3172\ : std_logic;
signal \N__3171\ : std_logic;
signal \N__3166\ : std_logic;
signal \N__3163\ : std_logic;
signal \N__3158\ : std_logic;
signal \N__3155\ : std_logic;
signal \N__3152\ : std_logic;
signal \N__3149\ : std_logic;
signal \N__3148\ : std_logic;
signal \N__3145\ : std_logic;
signal \N__3142\ : std_logic;
signal \N__3137\ : std_logic;
signal \N__3134\ : std_logic;
signal \N__3131\ : std_logic;
signal \N__3128\ : std_logic;
signal \N__3125\ : std_logic;
signal \N__3122\ : std_logic;
signal \N__3119\ : std_logic;
signal \N__3116\ : std_logic;
signal \N__3113\ : std_logic;
signal \N__3110\ : std_logic;
signal \N__3109\ : std_logic;
signal \N__3106\ : std_logic;
signal \N__3103\ : std_logic;
signal \N__3098\ : std_logic;
signal \N__3097\ : std_logic;
signal \N__3094\ : std_logic;
signal \N__3091\ : std_logic;
signal \N__3086\ : std_logic;
signal \N__3085\ : std_logic;
signal \N__3082\ : std_logic;
signal \N__3079\ : std_logic;
signal \N__3074\ : std_logic;
signal \N__3071\ : std_logic;
signal \N__3070\ : std_logic;
signal \N__3067\ : std_logic;
signal \N__3064\ : std_logic;
signal \N__3061\ : std_logic;
signal \N__3056\ : std_logic;
signal \N__3055\ : std_logic;
signal \N__3052\ : std_logic;
signal \N__3049\ : std_logic;
signal \N__3044\ : std_logic;
signal \N__3041\ : std_logic;
signal \N__3038\ : std_logic;
signal \N__3035\ : std_logic;
signal \N__3032\ : std_logic;
signal \N__3031\ : std_logic;
signal \N__3028\ : std_logic;
signal \N__3025\ : std_logic;
signal \N__3020\ : std_logic;
signal \N__3017\ : std_logic;
signal \N__3014\ : std_logic;
signal \N__3013\ : std_logic;
signal \N__3010\ : std_logic;
signal \N__3007\ : std_logic;
signal \N__3002\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2996\ : std_logic;
signal \N__2993\ : std_logic;
signal \N__2990\ : std_logic;
signal \N__2987\ : std_logic;
signal \N__2986\ : std_logic;
signal \N__2983\ : std_logic;
signal \N__2980\ : std_logic;
signal \N__2975\ : std_logic;
signal \N__2972\ : std_logic;
signal \N__2971\ : std_logic;
signal \N__2968\ : std_logic;
signal \N__2965\ : std_logic;
signal \N__2960\ : std_logic;
signal \N__2957\ : std_logic;
signal \N__2956\ : std_logic;
signal \N__2953\ : std_logic;
signal \N__2950\ : std_logic;
signal \N__2947\ : std_logic;
signal \N__2944\ : std_logic;
signal \N__2939\ : std_logic;
signal \N__2936\ : std_logic;
signal \N__2933\ : std_logic;
signal \N__2930\ : std_logic;
signal \N__2929\ : std_logic;
signal \N__2926\ : std_logic;
signal \N__2923\ : std_logic;
signal \N__2920\ : std_logic;
signal \N__2917\ : std_logic;
signal \N__2912\ : std_logic;
signal \N__2911\ : std_logic;
signal \N__2908\ : std_logic;
signal \N__2905\ : std_logic;
signal \N__2900\ : std_logic;
signal \N__2899\ : std_logic;
signal \N__2896\ : std_logic;
signal \N__2893\ : std_logic;
signal \N__2888\ : std_logic;
signal \N__2885\ : std_logic;
signal \N__2884\ : std_logic;
signal \N__2881\ : std_logic;
signal \N__2878\ : std_logic;
signal \N__2873\ : std_logic;
signal \N__2872\ : std_logic;
signal \N__2869\ : std_logic;
signal \N__2866\ : std_logic;
signal \N__2861\ : std_logic;
signal \N__2860\ : std_logic;
signal \N__2857\ : std_logic;
signal \N__2856\ : std_logic;
signal \N__2855\ : std_logic;
signal \N__2852\ : std_logic;
signal \N__2847\ : std_logic;
signal \N__2844\ : std_logic;
signal \N__2841\ : std_logic;
signal \N__2834\ : std_logic;
signal \N__2833\ : std_logic;
signal \N__2830\ : std_logic;
signal \N__2827\ : std_logic;
signal \N__2822\ : std_logic;
signal \N__2821\ : std_logic;
signal \N__2818\ : std_logic;
signal \N__2815\ : std_logic;
signal \N__2810\ : std_logic;
signal \N__2807\ : std_logic;
signal \N__2806\ : std_logic;
signal \N__2803\ : std_logic;
signal \N__2800\ : std_logic;
signal \N__2795\ : std_logic;
signal \N__2792\ : std_logic;
signal \N__2789\ : std_logic;
signal \N__2786\ : std_logic;
signal \N__2783\ : std_logic;
signal \N__2780\ : std_logic;
signal \N__2777\ : std_logic;
signal \N__2774\ : std_logic;
signal \N__2771\ : std_logic;
signal \N__2768\ : std_logic;
signal \N__2765\ : std_logic;
signal \N__2762\ : std_logic;
signal \N__2759\ : std_logic;
signal \N__2756\ : std_logic;
signal \N__2753\ : std_logic;
signal \N__2750\ : std_logic;
signal \N__2747\ : std_logic;
signal \N__2744\ : std_logic;
signal \N__2741\ : std_logic;
signal \N__2738\ : std_logic;
signal \N__2735\ : std_logic;
signal \N__2734\ : std_logic;
signal \N__2731\ : std_logic;
signal \N__2728\ : std_logic;
signal \N__2723\ : std_logic;
signal \N__2720\ : std_logic;
signal \N__2719\ : std_logic;
signal \N__2718\ : std_logic;
signal \N__2717\ : std_logic;
signal \N__2714\ : std_logic;
signal \N__2711\ : std_logic;
signal \N__2706\ : std_logic;
signal \N__2703\ : std_logic;
signal \N__2696\ : std_logic;
signal \N__2693\ : std_logic;
signal \N__2690\ : std_logic;
signal \N__2687\ : std_logic;
signal \N__2684\ : std_logic;
signal \N__2683\ : std_logic;
signal \N__2680\ : std_logic;
signal \N__2677\ : std_logic;
signal \N__2672\ : std_logic;
signal \N__2671\ : std_logic;
signal \N__2668\ : std_logic;
signal \N__2665\ : std_logic;
signal \N__2660\ : std_logic;
signal \N__2659\ : std_logic;
signal \N__2656\ : std_logic;
signal \N__2653\ : std_logic;
signal \N__2648\ : std_logic;
signal \N__2645\ : std_logic;
signal \N__2644\ : std_logic;
signal \N__2641\ : std_logic;
signal \N__2638\ : std_logic;
signal \N__2633\ : std_logic;
signal \N__2632\ : std_logic;
signal \N__2629\ : std_logic;
signal \N__2626\ : std_logic;
signal \N__2621\ : std_logic;
signal \N__2620\ : std_logic;
signal \N__2619\ : std_logic;
signal \N__2618\ : std_logic;
signal \N__2617\ : std_logic;
signal \N__2616\ : std_logic;
signal \N__2613\ : std_logic;
signal \N__2612\ : std_logic;
signal \N__2609\ : std_logic;
signal \N__2606\ : std_logic;
signal \N__2597\ : std_logic;
signal \N__2596\ : std_logic;
signal \N__2595\ : std_logic;
signal \N__2592\ : std_logic;
signal \N__2589\ : std_logic;
signal \N__2586\ : std_logic;
signal \N__2583\ : std_logic;
signal \N__2578\ : std_logic;
signal \N__2575\ : std_logic;
signal \N__2564\ : std_logic;
signal \N__2563\ : std_logic;
signal \N__2562\ : std_logic;
signal \N__2561\ : std_logic;
signal \N__2560\ : std_logic;
signal \N__2557\ : std_logic;
signal \N__2556\ : std_logic;
signal \N__2555\ : std_logic;
signal \N__2552\ : std_logic;
signal \N__2549\ : std_logic;
signal \N__2548\ : std_logic;
signal \N__2545\ : std_logic;
signal \N__2544\ : std_logic;
signal \N__2539\ : std_logic;
signal \N__2530\ : std_logic;
signal \N__2523\ : std_logic;
signal \N__2516\ : std_logic;
signal \N__2515\ : std_logic;
signal \N__2514\ : std_logic;
signal \N__2513\ : std_logic;
signal \N__2504\ : std_logic;
signal \N__2503\ : std_logic;
signal \N__2502\ : std_logic;
signal \N__2501\ : std_logic;
signal \N__2500\ : std_logic;
signal \N__2499\ : std_logic;
signal \N__2498\ : std_logic;
signal \N__2495\ : std_logic;
signal \N__2486\ : std_logic;
signal \N__2481\ : std_logic;
signal \N__2474\ : std_logic;
signal \N__2471\ : std_logic;
signal \N__2468\ : std_logic;
signal \N__2465\ : std_logic;
signal \N__2464\ : std_logic;
signal \N__2461\ : std_logic;
signal \N__2458\ : std_logic;
signal \N__2453\ : std_logic;
signal \N__2450\ : std_logic;
signal \N__2447\ : std_logic;
signal \N__2444\ : std_logic;
signal \N__2443\ : std_logic;
signal \N__2440\ : std_logic;
signal \N__2437\ : std_logic;
signal \N__2432\ : std_logic;
signal \N__2431\ : std_logic;
signal \N__2428\ : std_logic;
signal \N__2425\ : std_logic;
signal \N__2420\ : std_logic;
signal \N__2417\ : std_logic;
signal \N__2416\ : std_logic;
signal \N__2413\ : std_logic;
signal \N__2410\ : std_logic;
signal \N__2405\ : std_logic;
signal \N__2404\ : std_logic;
signal \N__2401\ : std_logic;
signal \N__2398\ : std_logic;
signal \N__2393\ : std_logic;
signal \N__2392\ : std_logic;
signal \N__2391\ : std_logic;
signal \N__2386\ : std_logic;
signal \N__2383\ : std_logic;
signal \N__2378\ : std_logic;
signal \N__2375\ : std_logic;
signal \N__2372\ : std_logic;
signal \N__2371\ : std_logic;
signal \N__2368\ : std_logic;
signal \N__2365\ : std_logic;
signal \N__2360\ : std_logic;
signal \N__2357\ : std_logic;
signal \N__2356\ : std_logic;
signal \N__2353\ : std_logic;
signal \N__2350\ : std_logic;
signal \N__2347\ : std_logic;
signal \N__2344\ : std_logic;
signal \N__2339\ : std_logic;
signal \N__2336\ : std_logic;
signal \N__2333\ : std_logic;
signal \N__2332\ : std_logic;
signal \N__2329\ : std_logic;
signal \N__2326\ : std_logic;
signal \N__2321\ : std_logic;
signal \N__2320\ : std_logic;
signal \N__2317\ : std_logic;
signal \N__2314\ : std_logic;
signal \N__2309\ : std_logic;
signal \N__2308\ : std_logic;
signal \N__2305\ : std_logic;
signal \N__2302\ : std_logic;
signal \N__2297\ : std_logic;
signal \N__2296\ : std_logic;
signal \N__2293\ : std_logic;
signal \N__2290\ : std_logic;
signal \N__2285\ : std_logic;
signal \N__2282\ : std_logic;
signal \N__2279\ : std_logic;
signal \N__2276\ : std_logic;
signal \N__2273\ : std_logic;
signal \N__2270\ : std_logic;
signal \N__2267\ : std_logic;
signal \N__2264\ : std_logic;
signal \N__2261\ : std_logic;
signal \N__2258\ : std_logic;
signal \N__2255\ : std_logic;
signal \N__2252\ : std_logic;
signal \N__2251\ : std_logic;
signal \N__2246\ : std_logic;
signal \N__2243\ : std_logic;
signal \N__2242\ : std_logic;
signal \N__2237\ : std_logic;
signal \N__2234\ : std_logic;
signal \N__2233\ : std_logic;
signal \N__2230\ : std_logic;
signal \N__2225\ : std_logic;
signal \N__2222\ : std_logic;
signal \N__2221\ : std_logic;
signal \N__2218\ : std_logic;
signal \N__2215\ : std_logic;
signal \N__2210\ : std_logic;
signal \N__2207\ : std_logic;
signal \N__2204\ : std_logic;
signal \N__2201\ : std_logic;
signal \N__2198\ : std_logic;
signal \N__2195\ : std_logic;
signal \N__2192\ : std_logic;
signal \N__2189\ : std_logic;
signal \N__2186\ : std_logic;
signal \N__2183\ : std_logic;
signal \N__2180\ : std_logic;
signal \N__2177\ : std_logic;
signal \N__2174\ : std_logic;
signal \N__2171\ : std_logic;
signal \N__2168\ : std_logic;
signal \N__2165\ : std_logic;
signal \N__2162\ : std_logic;
signal \N__2159\ : std_logic;
signal \N__2156\ : std_logic;
signal \N__2153\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \bfn_7_5_0_\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_5hz_cry_1\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_5hz_cry_2\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_5hz_cry_3\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_5hz_cry_4\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_5hz_cry_5\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_5hz_cry_6\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_5hz_cry_7\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_5hz_cry_8\ : std_logic;
signal \bfn_7_6_0_\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_5hz_cry_9\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_5hz_cry_10\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_5hz_cry_11\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_5hz_cry_12\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_5hz_cry_13\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_5hz_cry_14\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_5hz_cry_15\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_5hz_cry_16\ : std_logic;
signal \bfn_7_7_0_\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_5hz_cry_17\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_5hz_cry_18\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_5hz_cry_19\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_5hz_cry_20\ : std_logic;
signal \LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_18\ : std_logic;
signal \LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_21\ : std_logic;
signal \LED_Blink_Inst.r_Count_5HZZ0Z_19\ : std_logic;
signal \LED_Blink_Inst.r_Count_5HZZ0Z_20\ : std_logic;
signal \LED_Blink_Inst.r_Count_5HZZ0Z_21\ : std_logic;
signal \LED_Blink_Inst.r_Count_5HZZ0Z_15\ : std_logic;
signal \LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_7\ : std_logic;
signal \LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_5\ : std_logic;
signal \LED_Blink_Inst.r_Count_5HZZ0Z_4\ : std_logic;
signal \LED_Blink_Inst.r_Count_5HZZ0Z_2\ : std_logic;
signal \LED_Blink_Inst.r_Count_5HZZ0Z_6\ : std_logic;
signal \LED_Blink_Inst.r_Count_5HZZ0Z_7\ : std_logic;
signal \LED_Blink_Inst.r_Count_5HZZ0Z_1\ : std_logic;
signal \LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_8\ : std_logic;
signal \LED_Blink_Inst.r_Count_5HZZ0Z_8\ : std_logic;
signal \o_LED_2_c\ : std_logic;
signal \LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_13\ : std_logic;
signal \LED_Blink_Inst.r_Count_5HZZ0Z_13\ : std_logic;
signal \LED_Blink_Inst.r_Count_5HZZ0Z_18\ : std_logic;
signal \LED_Blink_Inst.r_Count_5HZZ0Z_5\ : std_logic;
signal \LED_Blink_Inst.r_Count_5HZZ0Z_3\ : std_logic;
signal \LED_Blink_Inst.un1_r_count_5hz_13_cascade_\ : std_logic;
signal \LED_Blink_Inst.un1_r_count_5hz_3\ : std_logic;
signal \LED_Blink_Inst.un1_r_count_5hz_11\ : std_logic;
signal \LED_Blink_Inst.r_Count_5HZZ0Z_11\ : std_logic;
signal \LED_Blink_Inst.un1_r_count_5hz_17_cascade_\ : std_logic;
signal \LED_Blink_Inst.r_Count_5HZZ0Z_0\ : std_logic;
signal \LED_Blink_Inst.un1_r_count_5hz_19_cascade_\ : std_logic;
signal \LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_17\ : std_logic;
signal \LED_Blink_Inst.r_Count_5HZZ0Z_17\ : std_logic;
signal \LED_Blink_Inst.r_Count_5HZZ0Z_9\ : std_logic;
signal \LED_Blink_Inst.r_Count_5HZZ0Z_14\ : std_logic;
signal \LED_Blink_Inst.r_Count_5HZZ0Z_16\ : std_logic;
signal \LED_Blink_Inst.r_Count_5HZZ0Z_12\ : std_logic;
signal \LED_Blink_Inst.un1_r_count_5hz_15\ : std_logic;
signal \LED_Blink_Inst.un1_r_count_5hz_19\ : std_logic;
signal \LED_Blink_Inst.un1_r_count_5hz_14\ : std_logic;
signal \LED_Blink_Inst.un1_r_count_5hz_15_cascade_\ : std_logic;
signal \LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_10\ : std_logic;
signal \LED_Blink_Inst.r_Count_5HZZ0Z_10\ : std_logic;
signal \bfn_8_7_0_\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_1hz_cry_1\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_1hz_cry_2\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_1hz_cry_3\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_1hz_cry_4\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_1hz_cry_5\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_1hz_cry_6\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_1hz_cry_7\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_1hz_cry_8\ : std_logic;
signal \bfn_8_8_0_\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_1hz_cry_9\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_1hz_cry_10\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_1hz_cry_11\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_1hz_cry_12\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_1hz_cry_13\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_1hz_cry_14\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_1hz_cry_15\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_1hz_cry_16\ : std_logic;
signal \bfn_8_9_0_\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_1hz_cry_17\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_1hz_cry_18\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_1hz_cry_19\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_1hz_cry_20\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_1hz_cry_21\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_1hz_cry_22\ : std_logic;
signal \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_23_cascade_\ : std_logic;
signal \LED_Blink_Inst.r_Count_1HZZ0Z_13\ : std_logic;
signal \LED_Blink_Inst.r_Count_1HZZ0Z_10\ : std_logic;
signal \LED_Blink_Inst.r_Count_1HZZ0Z_15\ : std_logic;
signal \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_8\ : std_logic;
signal \o_LED_4_c\ : std_logic;
signal \LED_Blink_Inst.r_Count_1HZZ0Z_5\ : std_logic;
signal \LED_Blink_Inst.r_Count_1HZZ0Z_6\ : std_logic;
signal \LED_Blink_Inst.r_Count_1HZZ0Z_7\ : std_logic;
signal \LED_Blink_Inst.r_Count_1HZZ0Z_4\ : std_logic;
signal \LED_Blink_Inst.r_Count_1HZZ0Z_0\ : std_logic;
signal \LED_Blink_Inst.r_Count_1HZZ0Z_3\ : std_logic;
signal \LED_Blink_Inst.r_Count_1HZZ0Z_2\ : std_logic;
signal \LED_Blink_Inst.r_Count_1HZZ0Z_8\ : std_logic;
signal \LED_Blink_Inst.r_Count_1HZZ0Z_1\ : std_logic;
signal \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_11\ : std_logic;
signal \LED_Blink_Inst.r_Count_1HZZ0Z_11\ : std_logic;
signal \LED_Blink_Inst.un1_r_count_1hz_13\ : std_logic;
signal \LED_Blink_Inst.un1_r_count_1hz_14_cascade_\ : std_logic;
signal \LED_Blink_Inst.un1_r_count_1hz_12\ : std_logic;
signal \LED_Blink_Inst.un1_r_count_1hz_21_cascade_\ : std_logic;
signal \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_12\ : std_logic;
signal \LED_Blink_Inst.r_Count_1HZZ0Z_12\ : std_logic;
signal \LED_Blink_Inst.r_Count_1HZZ0Z_22\ : std_logic;
signal \LED_Blink_Inst.r_Count_1HZZ0Z_19\ : std_logic;
signal \LED_Blink_Inst.r_Count_1HZZ0Z_23\ : std_logic;
signal \LED_Blink_Inst.r_Count_1HZZ0Z_14\ : std_logic;
signal \LED_Blink_Inst.un1_r_count_1hz_16_cascade_\ : std_logic;
signal \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_16\ : std_logic;
signal \LED_Blink_Inst.r_Count_1HZZ0Z_16\ : std_logic;
signal \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_9\ : std_logic;
signal \LED_Blink_Inst.r_Count_1HZZ0Z_9\ : std_logic;
signal \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_20\ : std_logic;
signal \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_18\ : std_logic;
signal \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_21\ : std_logic;
signal \LED_Blink_Inst.un1_r_count_1hz_21\ : std_logic;
signal \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_17\ : std_logic;
signal \LED_Blink_Inst.un1_r_count_1hz_17\ : std_logic;
signal \LED_Blink_Inst.un1_r_count_1hz_16\ : std_logic;
signal \LED_Blink_Inst.r_Count_1HZZ0Z_20\ : std_logic;
signal \LED_Blink_Inst.r_Count_1HZZ0Z_18\ : std_logic;
signal \LED_Blink_Inst.r_Count_1HZZ0Z_21\ : std_logic;
signal \LED_Blink_Inst.r_Count_1HZZ0Z_17\ : std_logic;
signal \LED_Blink_Inst.un1_r_count_1hz_15\ : std_logic;
signal \bfn_11_3_0_\ : std_logic;
signal \LED_Blink_Inst.un6_r_count_10hz_cry_1\ : std_logic;
signal \LED_Blink_Inst.un6_r_count_10hz_cry_2\ : std_logic;
signal \LED_Blink_Inst.un6_r_count_10hz_cry_3\ : std_logic;
signal \LED_Blink_Inst.un6_r_count_10hz_cry_4\ : std_logic;
signal \LED_Blink_Inst.un6_r_count_10hz_cry_5\ : std_logic;
signal \LED_Blink_Inst.un6_r_count_10hz_cry_6\ : std_logic;
signal \LED_Blink_Inst.un6_r_count_10hz_cry_7\ : std_logic;
signal \LED_Blink_Inst.un6_r_count_10hz_cry_8\ : std_logic;
signal \bfn_11_4_0_\ : std_logic;
signal \LED_Blink_Inst.un6_r_count_10hz_cry_9\ : std_logic;
signal \LED_Blink_Inst.un6_r_count_10hz_cry_10\ : std_logic;
signal \LED_Blink_Inst.un6_r_count_10hz_cry_11\ : std_logic;
signal \LED_Blink_Inst.un6_r_count_10hz_cry_12\ : std_logic;
signal \LED_Blink_Inst.un6_r_count_10hz_cry_13\ : std_logic;
signal \LED_Blink_Inst.un6_r_count_10hz_cry_14\ : std_logic;
signal \LED_Blink_Inst.un6_r_count_10hz_cry_15\ : std_logic;
signal \LED_Blink_Inst.un6_r_count_10hz_cry_16\ : std_logic;
signal \bfn_11_5_0_\ : std_logic;
signal \LED_Blink_Inst.un6_r_count_10hz_cry_17\ : std_logic;
signal \LED_Blink_Inst.un6_r_count_10hz_cry_18\ : std_logic;
signal \LED_Blink_Inst.un6_r_count_10hz_cry_19\ : std_logic;
signal \LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_20_cascade_\ : std_logic;
signal \LED_Blink_Inst.r_Count_10HZZ0Z_20\ : std_logic;
signal \LED_Blink_Inst.r_Count_10HZZ0Z_19\ : std_logic;
signal \LED_Blink_Inst.r_Count_10HZZ0Z_18\ : std_logic;
signal \LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_17\ : std_logic;
signal \LED_Blink_Inst.r_Count_10HZZ0Z_17\ : std_logic;
signal \LED_Blink_Inst.un1_r_count_2hz_11\ : std_logic;
signal \LED_Blink_Inst.un1_r_count_2hz_12\ : std_logic;
signal \LED_Blink_Inst.un1_r_count_2hz_14_cascade_\ : std_logic;
signal \LED_Blink_Inst.un1_r_count_2hz_13\ : std_logic;
signal \LED_Blink_Inst.un1_r_count_2hz_20_cascade_\ : std_logic;
signal \LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_7\ : std_logic;
signal \LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_4\ : std_logic;
signal \LED_Blink_Inst.r_Count_10HZZ0Z_5\ : std_logic;
signal \LED_Blink_Inst.r_Count_10HZZ0Z_3\ : std_logic;
signal \LED_Blink_Inst.r_Count_10HZZ0Z_0\ : std_logic;
signal \LED_Blink_Inst.r_Count_10HZZ0Z_4\ : std_logic;
signal \LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_6\ : std_logic;
signal \LED_Blink_Inst.r_Count_10HZZ0Z_6\ : std_logic;
signal \LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_16\ : std_logic;
signal \LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_12\ : std_logic;
signal \LED_Blink_Inst.r_Count_10HZZ0Z_13\ : std_logic;
signal \LED_Blink_Inst.r_Count_10HZZ0Z_15\ : std_logic;
signal \LED_Blink_Inst.r_Count_10HZZ0Z_14\ : std_logic;
signal \LED_Blink_Inst.r_Count_10HZZ0Z_11\ : std_logic;
signal \LED_Blink_Inst.r_Count_10HZZ0Z_12\ : std_logic;
signal \LED_Blink_Inst.r_Count_10HZZ0Z_7\ : std_logic;
signal \LED_Blink_Inst.r_Count_10HZZ0Z_16\ : std_logic;
signal \LED_Blink_Inst.r_Count_10HZZ0Z_2\ : std_logic;
signal \LED_Blink_Inst.r_Count_10HZZ0Z_1\ : std_logic;
signal \LED_Blink_Inst.un1_r_count_10hz_12_cascade_\ : std_logic;
signal \LED_Blink_Inst.un1_r_count_10hz_2\ : std_logic;
signal \LED_Blink_Inst.r_Count_10HZZ0Z_8\ : std_logic;
signal \LED_Blink_Inst.r_Count_10HZZ0Z_10\ : std_logic;
signal \LED_Blink_Inst.un1_r_count_10hz_16_cascade_\ : std_logic;
signal \LED_Blink_Inst.un1_r_count_10hz_10\ : std_logic;
signal \LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_9\ : std_logic;
signal \LED_Blink_Inst.un1_r_count_10hz_18_cascade_\ : std_logic;
signal \LED_Blink_Inst.r_Count_10HZZ0Z_9\ : std_logic;
signal \LED_Blink_Inst.un1_r_count_10hz_14\ : std_logic;
signal \LED_Blink_Inst.un1_r_count_10hz_13\ : std_logic;
signal \LED_Blink_Inst.un1_r_count_10hz_18\ : std_logic;
signal \o_LED_1_c\ : std_logic;
signal \LED_Blink_Inst.r_Count_2HZZ0Z_1\ : std_logic;
signal \LED_Blink_Inst.r_Count_2HZZ0Z_0\ : std_logic;
signal \bfn_12_6_0_\ : std_logic;
signal \LED_Blink_Inst.r_Count_2HZZ0Z_2\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_2hz_cry_1\ : std_logic;
signal \LED_Blink_Inst.r_Count_2HZZ0Z_3\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_2hz_cry_2\ : std_logic;
signal \LED_Blink_Inst.r_Count_2HZZ0Z_4\ : std_logic;
signal \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_4\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_2hz_cry_3\ : std_logic;
signal \LED_Blink_Inst.r_Count_2HZZ0Z_5\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_2hz_cry_4\ : std_logic;
signal \LED_Blink_Inst.r_Count_2HZZ0Z_6\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_2hz_cry_5\ : std_logic;
signal \LED_Blink_Inst.r_Count_2HZZ0Z_7\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_2hz_cry_6\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_2hz_cry_7\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_2hz_cry_8\ : std_logic;
signal \LED_Blink_Inst.r_Count_2HZZ0Z_9\ : std_logic;
signal \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_9\ : std_logic;
signal \bfn_12_7_0_\ : std_logic;
signal \LED_Blink_Inst.r_Count_2HZZ0Z_10\ : std_logic;
signal \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_10\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_2hz_cry_9\ : std_logic;
signal \LED_Blink_Inst.r_Count_2HZZ0Z_11\ : std_logic;
signal \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_11\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_2hz_cry_10\ : std_logic;
signal \LED_Blink_Inst.r_Count_2HZZ0Z_12\ : std_logic;
signal \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_12\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_2hz_cry_11\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_2hz_cry_12\ : std_logic;
signal \LED_Blink_Inst.r_Count_2HZZ0Z_14\ : std_logic;
signal \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_14\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_2hz_cry_13\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_2hz_cry_14\ : std_logic;
signal \LED_Blink_Inst.r_Count_2HZZ0Z_16\ : std_logic;
signal \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_16\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_2hz_cry_15\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_2hz_cry_16\ : std_logic;
signal \bfn_12_8_0_\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_2hz_cry_17\ : std_logic;
signal \LED_Blink_Inst.r_Count_2HZZ0Z_19\ : std_logic;
signal \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_19\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_2hz_cry_18\ : std_logic;
signal \LED_Blink_Inst.r_Count_2HZZ0Z_20\ : std_logic;
signal \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_20\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_2hz_cry_19\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_2hz_cry_20\ : std_logic;
signal \LED_Blink_Inst.un4_r_count_2hz_cry_21\ : std_logic;
signal \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_22_cascade_\ : std_logic;
signal \LED_Blink_Inst.r_Count_2HZZ0Z_22\ : std_logic;
signal \LED_Blink_Inst.r_Count_2HZZ0Z_15\ : std_logic;
signal \LED_Blink_Inst.r_Count_2HZZ0Z_13\ : std_logic;
signal \LED_Blink_Inst.r_Count_2HZZ0Z_21\ : std_logic;
signal \LED_Blink_Inst.r_Count_2HZZ0Z_8\ : std_logic;
signal \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_17\ : std_logic;
signal \LED_Blink_Inst.r_Count_2HZZ0Z_17\ : std_logic;
signal \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_18\ : std_logic;
signal \LED_Blink_Inst.r_Count_2HZZ0Z_18\ : std_logic;
signal \LED_Blink_Inst.un1_r_count_2hz_15\ : std_logic;
signal \LED_Blink_Inst.un1_r_count_2hz_16\ : std_logic;
signal \LED_Blink_Inst.un1_r_count_2hz_20\ : std_logic;
signal \o_LED_3_c\ : std_logic;
signal \i_Clk_c_g\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \i_Clk_wire\ : std_logic;
signal \o_LED_1_wire\ : std_logic;
signal \o_LED_2_wire\ : std_logic;
signal \o_LED_3_wire\ : std_logic;
signal \o_LED_4_wire\ : std_logic;

begin
    \i_Clk_wire\ <= i_Clk;
    o_LED_1 <= \o_LED_1_wire\;
    o_LED_2 <= \o_LED_2_wire\;
    o_LED_3 <= \o_LED_3_wire\;
    o_LED_4 <= \o_LED_4_wire\;

    \i_Clk_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__4821\,
            GLOBALBUFFEROUTPUT => \i_Clk_c_g\
        );

    \i_Clk_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4823\,
            DIN => \N__4822\,
            DOUT => \N__4821\,
            PACKAGEPIN => \i_Clk_wire\
        );

    \i_Clk_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4823\,
            PADOUT => \N__4822\,
            PADIN => \N__4821\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_LED_1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4812\,
            DIN => \N__4811\,
            DOUT => \N__4810\,
            PACKAGEPIN => \o_LED_1_wire\
        );

    \o_LED_1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4812\,
            PADOUT => \N__4811\,
            PADIN => \N__4810\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3796\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_LED_2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4803\,
            DIN => \N__4802\,
            DOUT => \N__4801\,
            PACKAGEPIN => \o_LED_2_wire\
        );

    \o_LED_2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4803\,
            PADOUT => \N__4802\,
            PADIN => \N__4801\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2360\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_LED_3_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4794\,
            DIN => \N__4793\,
            DOUT => \N__4792\,
            PACKAGEPIN => \o_LED_3_wire\
        );

    \o_LED_3_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4794\,
            PADOUT => \N__4793\,
            PADIN => \N__4792\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4466\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_LED_4_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4785\,
            DIN => \N__4784\,
            DOUT => \N__4783\,
            PACKAGEPIN => \o_LED_4_wire\
        );

    \o_LED_4_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4785\,
            PADOUT => \N__4784\,
            PADIN => \N__4783\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2933\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1055\ : InMux
    port map (
            O => \N__4766\,
            I => \LED_Blink_Inst.un4_r_count_2hz_cry_20\
        );

    \I__1054\ : InMux
    port map (
            O => \N__4763\,
            I => \LED_Blink_Inst.un4_r_count_2hz_cry_21\
        );

    \I__1053\ : CascadeMux
    port map (
            O => \N__4760\,
            I => \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_22_cascade_\
        );

    \I__1052\ : CascadeMux
    port map (
            O => \N__4757\,
            I => \N__4753\
        );

    \I__1051\ : InMux
    port map (
            O => \N__4756\,
            I => \N__4750\
        );

    \I__1050\ : InMux
    port map (
            O => \N__4753\,
            I => \N__4747\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__4750\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_22\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__4747\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_22\
        );

    \I__1047\ : InMux
    port map (
            O => \N__4742\,
            I => \N__4738\
        );

    \I__1046\ : InMux
    port map (
            O => \N__4741\,
            I => \N__4735\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__4738\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_15\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__4735\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_15\
        );

    \I__1043\ : InMux
    port map (
            O => \N__4730\,
            I => \N__4726\
        );

    \I__1042\ : InMux
    port map (
            O => \N__4729\,
            I => \N__4723\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__4726\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_13\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__4723\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_13\
        );

    \I__1039\ : CascadeMux
    port map (
            O => \N__4718\,
            I => \N__4715\
        );

    \I__1038\ : InMux
    port map (
            O => \N__4715\,
            I => \N__4709\
        );

    \I__1037\ : InMux
    port map (
            O => \N__4714\,
            I => \N__4709\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__4709\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_21\
        );

    \I__1035\ : InMux
    port map (
            O => \N__4706\,
            I => \N__4703\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__4703\,
            I => \N__4699\
        );

    \I__1033\ : InMux
    port map (
            O => \N__4702\,
            I => \N__4696\
        );

    \I__1032\ : Odrv4
    port map (
            O => \N__4699\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_8\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__4696\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_8\
        );

    \I__1030\ : CascadeMux
    port map (
            O => \N__4691\,
            I => \N__4688\
        );

    \I__1029\ : InMux
    port map (
            O => \N__4688\,
            I => \N__4685\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__4685\,
            I => \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_17\
        );

    \I__1027\ : CascadeMux
    port map (
            O => \N__4682\,
            I => \N__4679\
        );

    \I__1026\ : InMux
    port map (
            O => \N__4679\,
            I => \N__4675\
        );

    \I__1025\ : InMux
    port map (
            O => \N__4678\,
            I => \N__4672\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__4675\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_17\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__4672\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_17\
        );

    \I__1022\ : InMux
    port map (
            O => \N__4667\,
            I => \N__4664\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__4664\,
            I => \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_18\
        );

    \I__1020\ : InMux
    port map (
            O => \N__4661\,
            I => \N__4657\
        );

    \I__1019\ : InMux
    port map (
            O => \N__4660\,
            I => \N__4654\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__4657\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_18\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__4654\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_18\
        );

    \I__1016\ : InMux
    port map (
            O => \N__4649\,
            I => \N__4629\
        );

    \I__1015\ : InMux
    port map (
            O => \N__4648\,
            I => \N__4629\
        );

    \I__1014\ : InMux
    port map (
            O => \N__4647\,
            I => \N__4629\
        );

    \I__1013\ : InMux
    port map (
            O => \N__4646\,
            I => \N__4626\
        );

    \I__1012\ : InMux
    port map (
            O => \N__4645\,
            I => \N__4617\
        );

    \I__1011\ : InMux
    port map (
            O => \N__4644\,
            I => \N__4617\
        );

    \I__1010\ : InMux
    port map (
            O => \N__4643\,
            I => \N__4617\
        );

    \I__1009\ : InMux
    port map (
            O => \N__4642\,
            I => \N__4617\
        );

    \I__1008\ : InMux
    port map (
            O => \N__4641\,
            I => \N__4614\
        );

    \I__1007\ : InMux
    port map (
            O => \N__4640\,
            I => \N__4603\
        );

    \I__1006\ : InMux
    port map (
            O => \N__4639\,
            I => \N__4603\
        );

    \I__1005\ : InMux
    port map (
            O => \N__4638\,
            I => \N__4603\
        );

    \I__1004\ : InMux
    port map (
            O => \N__4637\,
            I => \N__4603\
        );

    \I__1003\ : InMux
    port map (
            O => \N__4636\,
            I => \N__4603\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__4629\,
            I => \LED_Blink_Inst.un1_r_count_2hz_15\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__4626\,
            I => \LED_Blink_Inst.un1_r_count_2hz_15\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__4617\,
            I => \LED_Blink_Inst.un1_r_count_2hz_15\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__4614\,
            I => \LED_Blink_Inst.un1_r_count_2hz_15\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__4603\,
            I => \LED_Blink_Inst.un1_r_count_2hz_15\
        );

    \I__997\ : CascadeMux
    port map (
            O => \N__4592\,
            I => \N__4587\
        );

    \I__996\ : CascadeMux
    port map (
            O => \N__4591\,
            I => \N__4581\
        );

    \I__995\ : CascadeMux
    port map (
            O => \N__4590\,
            I => \N__4575\
        );

    \I__994\ : InMux
    port map (
            O => \N__4587\,
            I => \N__4563\
        );

    \I__993\ : InMux
    port map (
            O => \N__4586\,
            I => \N__4563\
        );

    \I__992\ : InMux
    port map (
            O => \N__4585\,
            I => \N__4563\
        );

    \I__991\ : InMux
    port map (
            O => \N__4584\,
            I => \N__4552\
        );

    \I__990\ : InMux
    port map (
            O => \N__4581\,
            I => \N__4552\
        );

    \I__989\ : InMux
    port map (
            O => \N__4580\,
            I => \N__4552\
        );

    \I__988\ : InMux
    port map (
            O => \N__4579\,
            I => \N__4552\
        );

    \I__987\ : InMux
    port map (
            O => \N__4578\,
            I => \N__4552\
        );

    \I__986\ : InMux
    port map (
            O => \N__4575\,
            I => \N__4541\
        );

    \I__985\ : InMux
    port map (
            O => \N__4574\,
            I => \N__4541\
        );

    \I__984\ : InMux
    port map (
            O => \N__4573\,
            I => \N__4541\
        );

    \I__983\ : InMux
    port map (
            O => \N__4572\,
            I => \N__4541\
        );

    \I__982\ : InMux
    port map (
            O => \N__4571\,
            I => \N__4541\
        );

    \I__981\ : InMux
    port map (
            O => \N__4570\,
            I => \N__4538\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__4563\,
            I => \LED_Blink_Inst.un1_r_count_2hz_16\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__4552\,
            I => \LED_Blink_Inst.un1_r_count_2hz_16\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__4541\,
            I => \LED_Blink_Inst.un1_r_count_2hz_16\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__4538\,
            I => \LED_Blink_Inst.un1_r_count_2hz_16\
        );

    \I__976\ : CascadeMux
    port map (
            O => \N__4529\,
            I => \N__4525\
        );

    \I__975\ : CascadeMux
    port map (
            O => \N__4528\,
            I => \N__4521\
        );

    \I__974\ : InMux
    port map (
            O => \N__4525\,
            I => \N__4506\
        );

    \I__973\ : InMux
    port map (
            O => \N__4524\,
            I => \N__4506\
        );

    \I__972\ : InMux
    port map (
            O => \N__4521\,
            I => \N__4499\
        );

    \I__971\ : InMux
    port map (
            O => \N__4520\,
            I => \N__4499\
        );

    \I__970\ : InMux
    port map (
            O => \N__4519\,
            I => \N__4499\
        );

    \I__969\ : InMux
    port map (
            O => \N__4518\,
            I => \N__4496\
        );

    \I__968\ : InMux
    port map (
            O => \N__4517\,
            I => \N__4489\
        );

    \I__967\ : InMux
    port map (
            O => \N__4516\,
            I => \N__4489\
        );

    \I__966\ : InMux
    port map (
            O => \N__4515\,
            I => \N__4489\
        );

    \I__965\ : InMux
    port map (
            O => \N__4514\,
            I => \N__4480\
        );

    \I__964\ : InMux
    port map (
            O => \N__4513\,
            I => \N__4480\
        );

    \I__963\ : InMux
    port map (
            O => \N__4512\,
            I => \N__4480\
        );

    \I__962\ : InMux
    port map (
            O => \N__4511\,
            I => \N__4480\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__4506\,
            I => \N__4475\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__4499\,
            I => \N__4475\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__4496\,
            I => \LED_Blink_Inst.un1_r_count_2hz_20\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__4489\,
            I => \LED_Blink_Inst.un1_r_count_2hz_20\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__4480\,
            I => \LED_Blink_Inst.un1_r_count_2hz_20\
        );

    \I__956\ : Odrv4
    port map (
            O => \N__4475\,
            I => \LED_Blink_Inst.un1_r_count_2hz_20\
        );

    \I__955\ : IoInMux
    port map (
            O => \N__4466\,
            I => \N__4463\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__4463\,
            I => \N__4459\
        );

    \I__953\ : CascadeMux
    port map (
            O => \N__4462\,
            I => \N__4456\
        );

    \I__952\ : Span4Mux_s0_h
    port map (
            O => \N__4459\,
            I => \N__4453\
        );

    \I__951\ : InMux
    port map (
            O => \N__4456\,
            I => \N__4450\
        );

    \I__950\ : Odrv4
    port map (
            O => \N__4453\,
            I => \o_LED_3_c\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__4450\,
            I => \o_LED_3_c\
        );

    \I__948\ : ClkMux
    port map (
            O => \N__4445\,
            I => \N__4373\
        );

    \I__947\ : ClkMux
    port map (
            O => \N__4444\,
            I => \N__4373\
        );

    \I__946\ : ClkMux
    port map (
            O => \N__4443\,
            I => \N__4373\
        );

    \I__945\ : ClkMux
    port map (
            O => \N__4442\,
            I => \N__4373\
        );

    \I__944\ : ClkMux
    port map (
            O => \N__4441\,
            I => \N__4373\
        );

    \I__943\ : ClkMux
    port map (
            O => \N__4440\,
            I => \N__4373\
        );

    \I__942\ : ClkMux
    port map (
            O => \N__4439\,
            I => \N__4373\
        );

    \I__941\ : ClkMux
    port map (
            O => \N__4438\,
            I => \N__4373\
        );

    \I__940\ : ClkMux
    port map (
            O => \N__4437\,
            I => \N__4373\
        );

    \I__939\ : ClkMux
    port map (
            O => \N__4436\,
            I => \N__4373\
        );

    \I__938\ : ClkMux
    port map (
            O => \N__4435\,
            I => \N__4373\
        );

    \I__937\ : ClkMux
    port map (
            O => \N__4434\,
            I => \N__4373\
        );

    \I__936\ : ClkMux
    port map (
            O => \N__4433\,
            I => \N__4373\
        );

    \I__935\ : ClkMux
    port map (
            O => \N__4432\,
            I => \N__4373\
        );

    \I__934\ : ClkMux
    port map (
            O => \N__4431\,
            I => \N__4373\
        );

    \I__933\ : ClkMux
    port map (
            O => \N__4430\,
            I => \N__4373\
        );

    \I__932\ : ClkMux
    port map (
            O => \N__4429\,
            I => \N__4373\
        );

    \I__931\ : ClkMux
    port map (
            O => \N__4428\,
            I => \N__4373\
        );

    \I__930\ : ClkMux
    port map (
            O => \N__4427\,
            I => \N__4373\
        );

    \I__929\ : ClkMux
    port map (
            O => \N__4426\,
            I => \N__4373\
        );

    \I__928\ : ClkMux
    port map (
            O => \N__4425\,
            I => \N__4373\
        );

    \I__927\ : ClkMux
    port map (
            O => \N__4424\,
            I => \N__4373\
        );

    \I__926\ : ClkMux
    port map (
            O => \N__4423\,
            I => \N__4373\
        );

    \I__925\ : ClkMux
    port map (
            O => \N__4422\,
            I => \N__4373\
        );

    \I__924\ : GlobalMux
    port map (
            O => \N__4373\,
            I => \N__4370\
        );

    \I__923\ : gio2CtrlBuf
    port map (
            O => \N__4370\,
            I => \i_Clk_c_g\
        );

    \I__922\ : InMux
    port map (
            O => \N__4367\,
            I => \N__4363\
        );

    \I__921\ : InMux
    port map (
            O => \N__4366\,
            I => \N__4360\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__4363\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_12\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__4360\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_12\
        );

    \I__918\ : CascadeMux
    port map (
            O => \N__4355\,
            I => \N__4352\
        );

    \I__917\ : InMux
    port map (
            O => \N__4352\,
            I => \N__4349\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__4349\,
            I => \N__4346\
        );

    \I__915\ : Span4Mux_v
    port map (
            O => \N__4346\,
            I => \N__4343\
        );

    \I__914\ : Odrv4
    port map (
            O => \N__4343\,
            I => \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_12\
        );

    \I__913\ : InMux
    port map (
            O => \N__4340\,
            I => \LED_Blink_Inst.un4_r_count_2hz_cry_11\
        );

    \I__912\ : InMux
    port map (
            O => \N__4337\,
            I => \LED_Blink_Inst.un4_r_count_2hz_cry_12\
        );

    \I__911\ : InMux
    port map (
            O => \N__4334\,
            I => \N__4330\
        );

    \I__910\ : InMux
    port map (
            O => \N__4333\,
            I => \N__4327\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__4330\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_14\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__4327\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_14\
        );

    \I__907\ : InMux
    port map (
            O => \N__4322\,
            I => \N__4319\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__4319\,
            I => \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_14\
        );

    \I__905\ : InMux
    port map (
            O => \N__4316\,
            I => \LED_Blink_Inst.un4_r_count_2hz_cry_13\
        );

    \I__904\ : InMux
    port map (
            O => \N__4313\,
            I => \LED_Blink_Inst.un4_r_count_2hz_cry_14\
        );

    \I__903\ : InMux
    port map (
            O => \N__4310\,
            I => \N__4306\
        );

    \I__902\ : InMux
    port map (
            O => \N__4309\,
            I => \N__4303\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__4306\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_16\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__4303\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_16\
        );

    \I__899\ : CascadeMux
    port map (
            O => \N__4298\,
            I => \N__4295\
        );

    \I__898\ : InMux
    port map (
            O => \N__4295\,
            I => \N__4292\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__4292\,
            I => \N__4289\
        );

    \I__896\ : Odrv4
    port map (
            O => \N__4289\,
            I => \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_16\
        );

    \I__895\ : InMux
    port map (
            O => \N__4286\,
            I => \LED_Blink_Inst.un4_r_count_2hz_cry_15\
        );

    \I__894\ : InMux
    port map (
            O => \N__4283\,
            I => \bfn_12_8_0_\
        );

    \I__893\ : InMux
    port map (
            O => \N__4280\,
            I => \LED_Blink_Inst.un4_r_count_2hz_cry_17\
        );

    \I__892\ : InMux
    port map (
            O => \N__4277\,
            I => \N__4273\
        );

    \I__891\ : InMux
    port map (
            O => \N__4276\,
            I => \N__4270\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__4273\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_19\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__4270\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_19\
        );

    \I__888\ : CascadeMux
    port map (
            O => \N__4265\,
            I => \N__4262\
        );

    \I__887\ : InMux
    port map (
            O => \N__4262\,
            I => \N__4259\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__4259\,
            I => \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_19\
        );

    \I__885\ : InMux
    port map (
            O => \N__4256\,
            I => \LED_Blink_Inst.un4_r_count_2hz_cry_18\
        );

    \I__884\ : InMux
    port map (
            O => \N__4253\,
            I => \N__4249\
        );

    \I__883\ : InMux
    port map (
            O => \N__4252\,
            I => \N__4246\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__4249\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_20\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__4246\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_20\
        );

    \I__880\ : InMux
    port map (
            O => \N__4241\,
            I => \N__4238\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__4238\,
            I => \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_20\
        );

    \I__878\ : InMux
    port map (
            O => \N__4235\,
            I => \LED_Blink_Inst.un4_r_count_2hz_cry_19\
        );

    \I__877\ : InMux
    port map (
            O => \N__4232\,
            I => \N__4228\
        );

    \I__876\ : InMux
    port map (
            O => \N__4231\,
            I => \N__4225\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__4228\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_4\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__4225\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_4\
        );

    \I__873\ : CascadeMux
    port map (
            O => \N__4220\,
            I => \N__4217\
        );

    \I__872\ : InMux
    port map (
            O => \N__4217\,
            I => \N__4214\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__4214\,
            I => \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_4\
        );

    \I__870\ : InMux
    port map (
            O => \N__4211\,
            I => \LED_Blink_Inst.un4_r_count_2hz_cry_3\
        );

    \I__869\ : CascadeMux
    port map (
            O => \N__4208\,
            I => \N__4205\
        );

    \I__868\ : InMux
    port map (
            O => \N__4205\,
            I => \N__4201\
        );

    \I__867\ : InMux
    port map (
            O => \N__4204\,
            I => \N__4198\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__4201\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_5\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__4198\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_5\
        );

    \I__864\ : InMux
    port map (
            O => \N__4193\,
            I => \LED_Blink_Inst.un4_r_count_2hz_cry_4\
        );

    \I__863\ : InMux
    port map (
            O => \N__4190\,
            I => \N__4186\
        );

    \I__862\ : InMux
    port map (
            O => \N__4189\,
            I => \N__4183\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__4186\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_6\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__4183\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_6\
        );

    \I__859\ : InMux
    port map (
            O => \N__4178\,
            I => \LED_Blink_Inst.un4_r_count_2hz_cry_5\
        );

    \I__858\ : InMux
    port map (
            O => \N__4175\,
            I => \N__4171\
        );

    \I__857\ : InMux
    port map (
            O => \N__4174\,
            I => \N__4168\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__4171\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_7\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__4168\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_7\
        );

    \I__854\ : InMux
    port map (
            O => \N__4163\,
            I => \LED_Blink_Inst.un4_r_count_2hz_cry_6\
        );

    \I__853\ : InMux
    port map (
            O => \N__4160\,
            I => \LED_Blink_Inst.un4_r_count_2hz_cry_7\
        );

    \I__852\ : InMux
    port map (
            O => \N__4157\,
            I => \N__4153\
        );

    \I__851\ : InMux
    port map (
            O => \N__4156\,
            I => \N__4150\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__4153\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_9\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__4150\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_9\
        );

    \I__848\ : InMux
    port map (
            O => \N__4145\,
            I => \N__4142\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__4142\,
            I => \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_9\
        );

    \I__846\ : InMux
    port map (
            O => \N__4139\,
            I => \bfn_12_7_0_\
        );

    \I__845\ : InMux
    port map (
            O => \N__4136\,
            I => \N__4132\
        );

    \I__844\ : InMux
    port map (
            O => \N__4135\,
            I => \N__4129\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__4132\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_10\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__4129\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_10\
        );

    \I__841\ : CascadeMux
    port map (
            O => \N__4124\,
            I => \N__4121\
        );

    \I__840\ : InMux
    port map (
            O => \N__4121\,
            I => \N__4118\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__4118\,
            I => \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_10\
        );

    \I__838\ : InMux
    port map (
            O => \N__4115\,
            I => \LED_Blink_Inst.un4_r_count_2hz_cry_9\
        );

    \I__837\ : CascadeMux
    port map (
            O => \N__4112\,
            I => \N__4109\
        );

    \I__836\ : InMux
    port map (
            O => \N__4109\,
            I => \N__4105\
        );

    \I__835\ : InMux
    port map (
            O => \N__4108\,
            I => \N__4102\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__4105\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_11\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__4102\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_11\
        );

    \I__832\ : InMux
    port map (
            O => \N__4097\,
            I => \N__4094\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__4094\,
            I => \N__4091\
        );

    \I__830\ : Odrv4
    port map (
            O => \N__4091\,
            I => \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_11\
        );

    \I__829\ : InMux
    port map (
            O => \N__4088\,
            I => \LED_Blink_Inst.un4_r_count_2hz_cry_10\
        );

    \I__828\ : InMux
    port map (
            O => \N__4085\,
            I => \N__4081\
        );

    \I__827\ : InMux
    port map (
            O => \N__4084\,
            I => \N__4078\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__4081\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_12\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__4078\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_12\
        );

    \I__824\ : CascadeMux
    port map (
            O => \N__4073\,
            I => \N__4069\
        );

    \I__823\ : InMux
    port map (
            O => \N__4072\,
            I => \N__4066\
        );

    \I__822\ : InMux
    port map (
            O => \N__4069\,
            I => \N__4063\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__4066\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_7\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__4063\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_7\
        );

    \I__819\ : InMux
    port map (
            O => \N__4058\,
            I => \N__4054\
        );

    \I__818\ : InMux
    port map (
            O => \N__4057\,
            I => \N__4051\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__4054\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_16\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__4051\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_16\
        );

    \I__815\ : InMux
    port map (
            O => \N__4046\,
            I => \N__4042\
        );

    \I__814\ : InMux
    port map (
            O => \N__4045\,
            I => \N__4039\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__4042\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_2\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__4039\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_2\
        );

    \I__811\ : InMux
    port map (
            O => \N__4034\,
            I => \N__4029\
        );

    \I__810\ : InMux
    port map (
            O => \N__4033\,
            I => \N__4026\
        );

    \I__809\ : InMux
    port map (
            O => \N__4032\,
            I => \N__4023\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__4029\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_1\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__4026\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_1\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__4023\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_1\
        );

    \I__805\ : CascadeMux
    port map (
            O => \N__4016\,
            I => \LED_Blink_Inst.un1_r_count_10hz_12_cascade_\
        );

    \I__804\ : InMux
    port map (
            O => \N__4013\,
            I => \N__4010\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__4010\,
            I => \LED_Blink_Inst.un1_r_count_10hz_2\
        );

    \I__802\ : InMux
    port map (
            O => \N__4007\,
            I => \N__4003\
        );

    \I__801\ : InMux
    port map (
            O => \N__4006\,
            I => \N__4000\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__4003\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_8\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__4000\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_8\
        );

    \I__798\ : InMux
    port map (
            O => \N__3995\,
            I => \N__3991\
        );

    \I__797\ : InMux
    port map (
            O => \N__3994\,
            I => \N__3988\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__3991\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_10\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__3988\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_10\
        );

    \I__794\ : CascadeMux
    port map (
            O => \N__3983\,
            I => \LED_Blink_Inst.un1_r_count_10hz_16_cascade_\
        );

    \I__793\ : InMux
    port map (
            O => \N__3980\,
            I => \N__3977\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__3977\,
            I => \N__3974\
        );

    \I__791\ : Odrv4
    port map (
            O => \N__3974\,
            I => \LED_Blink_Inst.un1_r_count_10hz_10\
        );

    \I__790\ : InMux
    port map (
            O => \N__3971\,
            I => \N__3968\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__3968\,
            I => \LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_9\
        );

    \I__788\ : CascadeMux
    port map (
            O => \N__3965\,
            I => \LED_Blink_Inst.un1_r_count_10hz_18_cascade_\
        );

    \I__787\ : InMux
    port map (
            O => \N__3962\,
            I => \N__3958\
        );

    \I__786\ : InMux
    port map (
            O => \N__3961\,
            I => \N__3955\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__3958\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_9\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__3955\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_9\
        );

    \I__783\ : CascadeMux
    port map (
            O => \N__3950\,
            I => \N__3942\
        );

    \I__782\ : CascadeMux
    port map (
            O => \N__3949\,
            I => \N__3936\
        );

    \I__781\ : CascadeMux
    port map (
            O => \N__3948\,
            I => \N__3933\
        );

    \I__780\ : CascadeMux
    port map (
            O => \N__3947\,
            I => \N__3929\
        );

    \I__779\ : CascadeMux
    port map (
            O => \N__3946\,
            I => \N__3926\
        );

    \I__778\ : InMux
    port map (
            O => \N__3945\,
            I => \N__3921\
        );

    \I__777\ : InMux
    port map (
            O => \N__3942\,
            I => \N__3921\
        );

    \I__776\ : InMux
    port map (
            O => \N__3941\,
            I => \N__3918\
        );

    \I__775\ : InMux
    port map (
            O => \N__3940\,
            I => \N__3909\
        );

    \I__774\ : InMux
    port map (
            O => \N__3939\,
            I => \N__3909\
        );

    \I__773\ : InMux
    port map (
            O => \N__3936\,
            I => \N__3909\
        );

    \I__772\ : InMux
    port map (
            O => \N__3933\,
            I => \N__3909\
        );

    \I__771\ : InMux
    port map (
            O => \N__3932\,
            I => \N__3902\
        );

    \I__770\ : InMux
    port map (
            O => \N__3929\,
            I => \N__3902\
        );

    \I__769\ : InMux
    port map (
            O => \N__3926\,
            I => \N__3902\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__3921\,
            I => \LED_Blink_Inst.un1_r_count_10hz_14\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__3918\,
            I => \LED_Blink_Inst.un1_r_count_10hz_14\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__3909\,
            I => \LED_Blink_Inst.un1_r_count_10hz_14\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__3902\,
            I => \LED_Blink_Inst.un1_r_count_10hz_14\
        );

    \I__764\ : CascadeMux
    port map (
            O => \N__3893\,
            I => \N__3889\
        );

    \I__763\ : CascadeMux
    port map (
            O => \N__3892\,
            I => \N__3886\
        );

    \I__762\ : InMux
    port map (
            O => \N__3889\,
            I => \N__3871\
        );

    \I__761\ : InMux
    port map (
            O => \N__3886\,
            I => \N__3871\
        );

    \I__760\ : InMux
    port map (
            O => \N__3885\,
            I => \N__3871\
        );

    \I__759\ : InMux
    port map (
            O => \N__3884\,
            I => \N__3868\
        );

    \I__758\ : InMux
    port map (
            O => \N__3883\,
            I => \N__3865\
        );

    \I__757\ : InMux
    port map (
            O => \N__3882\,
            I => \N__3862\
        );

    \I__756\ : InMux
    port map (
            O => \N__3881\,
            I => \N__3857\
        );

    \I__755\ : InMux
    port map (
            O => \N__3880\,
            I => \N__3857\
        );

    \I__754\ : InMux
    port map (
            O => \N__3879\,
            I => \N__3852\
        );

    \I__753\ : InMux
    port map (
            O => \N__3878\,
            I => \N__3852\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__3871\,
            I => \N__3847\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__3868\,
            I => \N__3847\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__3865\,
            I => \LED_Blink_Inst.un1_r_count_10hz_13\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__3862\,
            I => \LED_Blink_Inst.un1_r_count_10hz_13\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__3857\,
            I => \LED_Blink_Inst.un1_r_count_10hz_13\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__3852\,
            I => \LED_Blink_Inst.un1_r_count_10hz_13\
        );

    \I__746\ : Odrv4
    port map (
            O => \N__3847\,
            I => \LED_Blink_Inst.un1_r_count_10hz_13\
        );

    \I__745\ : InMux
    port map (
            O => \N__3836\,
            I => \N__3825\
        );

    \I__744\ : InMux
    port map (
            O => \N__3835\,
            I => \N__3820\
        );

    \I__743\ : InMux
    port map (
            O => \N__3834\,
            I => \N__3820\
        );

    \I__742\ : InMux
    port map (
            O => \N__3833\,
            I => \N__3815\
        );

    \I__741\ : InMux
    port map (
            O => \N__3832\,
            I => \N__3815\
        );

    \I__740\ : InMux
    port map (
            O => \N__3831\,
            I => \N__3806\
        );

    \I__739\ : InMux
    port map (
            O => \N__3830\,
            I => \N__3806\
        );

    \I__738\ : InMux
    port map (
            O => \N__3829\,
            I => \N__3806\
        );

    \I__737\ : InMux
    port map (
            O => \N__3828\,
            I => \N__3806\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__3825\,
            I => \LED_Blink_Inst.un1_r_count_10hz_18\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__3820\,
            I => \LED_Blink_Inst.un1_r_count_10hz_18\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__3815\,
            I => \LED_Blink_Inst.un1_r_count_10hz_18\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__3806\,
            I => \LED_Blink_Inst.un1_r_count_10hz_18\
        );

    \I__732\ : CascadeMux
    port map (
            O => \N__3797\,
            I => \N__3793\
        );

    \I__731\ : IoInMux
    port map (
            O => \N__3796\,
            I => \N__3790\
        );

    \I__730\ : InMux
    port map (
            O => \N__3793\,
            I => \N__3787\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__3790\,
            I => \o_LED_1_c\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__3787\,
            I => \o_LED_1_c\
        );

    \I__727\ : InMux
    port map (
            O => \N__3782\,
            I => \N__3777\
        );

    \I__726\ : InMux
    port map (
            O => \N__3781\,
            I => \N__3774\
        );

    \I__725\ : InMux
    port map (
            O => \N__3780\,
            I => \N__3771\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__3777\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_1\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__3774\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_1\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__3771\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_1\
        );

    \I__721\ : CascadeMux
    port map (
            O => \N__3764\,
            I => \N__3758\
        );

    \I__720\ : InMux
    port map (
            O => \N__3763\,
            I => \N__3755\
        );

    \I__719\ : InMux
    port map (
            O => \N__3762\,
            I => \N__3750\
        );

    \I__718\ : InMux
    port map (
            O => \N__3761\,
            I => \N__3750\
        );

    \I__717\ : InMux
    port map (
            O => \N__3758\,
            I => \N__3747\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__3755\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_0\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__3750\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_0\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__3747\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_0\
        );

    \I__713\ : InMux
    port map (
            O => \N__3740\,
            I => \N__3736\
        );

    \I__712\ : InMux
    port map (
            O => \N__3739\,
            I => \N__3733\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__3736\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_2\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__3733\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_2\
        );

    \I__709\ : InMux
    port map (
            O => \N__3728\,
            I => \LED_Blink_Inst.un4_r_count_2hz_cry_1\
        );

    \I__708\ : InMux
    port map (
            O => \N__3725\,
            I => \N__3721\
        );

    \I__707\ : InMux
    port map (
            O => \N__3724\,
            I => \N__3718\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__3721\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_3\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__3718\,
            I => \LED_Blink_Inst.r_Count_2HZZ0Z_3\
        );

    \I__704\ : InMux
    port map (
            O => \N__3713\,
            I => \LED_Blink_Inst.un4_r_count_2hz_cry_2\
        );

    \I__703\ : InMux
    port map (
            O => \N__3710\,
            I => \N__3707\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__3707\,
            I => \LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_4\
        );

    \I__701\ : InMux
    port map (
            O => \N__3704\,
            I => \N__3700\
        );

    \I__700\ : InMux
    port map (
            O => \N__3703\,
            I => \N__3697\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__3700\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_5\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__3697\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_5\
        );

    \I__697\ : InMux
    port map (
            O => \N__3692\,
            I => \N__3688\
        );

    \I__696\ : InMux
    port map (
            O => \N__3691\,
            I => \N__3685\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__3688\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_3\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__3685\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_3\
        );

    \I__693\ : CascadeMux
    port map (
            O => \N__3680\,
            I => \N__3674\
        );

    \I__692\ : InMux
    port map (
            O => \N__3679\,
            I => \N__3667\
        );

    \I__691\ : InMux
    port map (
            O => \N__3678\,
            I => \N__3667\
        );

    \I__690\ : InMux
    port map (
            O => \N__3677\,
            I => \N__3667\
        );

    \I__689\ : InMux
    port map (
            O => \N__3674\,
            I => \N__3664\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__3667\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_0\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__3664\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_0\
        );

    \I__686\ : InMux
    port map (
            O => \N__3659\,
            I => \N__3655\
        );

    \I__685\ : InMux
    port map (
            O => \N__3658\,
            I => \N__3652\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__3655\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_4\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__3652\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_4\
        );

    \I__682\ : InMux
    port map (
            O => \N__3647\,
            I => \N__3644\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__3644\,
            I => \LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_6\
        );

    \I__680\ : InMux
    port map (
            O => \N__3641\,
            I => \N__3637\
        );

    \I__679\ : InMux
    port map (
            O => \N__3640\,
            I => \N__3634\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__3637\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_6\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__3634\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_6\
        );

    \I__676\ : InMux
    port map (
            O => \N__3629\,
            I => \N__3626\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__3626\,
            I => \LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_16\
        );

    \I__674\ : InMux
    port map (
            O => \N__3623\,
            I => \N__3620\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__3620\,
            I => \LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_12\
        );

    \I__672\ : InMux
    port map (
            O => \N__3617\,
            I => \N__3613\
        );

    \I__671\ : InMux
    port map (
            O => \N__3616\,
            I => \N__3610\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__3613\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_13\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__3610\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_13\
        );

    \I__668\ : InMux
    port map (
            O => \N__3605\,
            I => \N__3601\
        );

    \I__667\ : InMux
    port map (
            O => \N__3604\,
            I => \N__3598\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__3601\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_15\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__3598\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_15\
        );

    \I__664\ : CascadeMux
    port map (
            O => \N__3593\,
            I => \N__3590\
        );

    \I__663\ : InMux
    port map (
            O => \N__3590\,
            I => \N__3586\
        );

    \I__662\ : InMux
    port map (
            O => \N__3589\,
            I => \N__3583\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__3586\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_14\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__3583\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_14\
        );

    \I__659\ : InMux
    port map (
            O => \N__3578\,
            I => \N__3574\
        );

    \I__658\ : InMux
    port map (
            O => \N__3577\,
            I => \N__3571\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__3574\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_11\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__3571\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_11\
        );

    \I__655\ : InMux
    port map (
            O => \N__3566\,
            I => \N__3563\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__3563\,
            I => \LED_Blink_Inst.un1_r_count_2hz_11\
        );

    \I__653\ : InMux
    port map (
            O => \N__3560\,
            I => \N__3557\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__3557\,
            I => \LED_Blink_Inst.un1_r_count_2hz_12\
        );

    \I__651\ : CascadeMux
    port map (
            O => \N__3554\,
            I => \LED_Blink_Inst.un1_r_count_2hz_14_cascade_\
        );

    \I__650\ : InMux
    port map (
            O => \N__3551\,
            I => \N__3548\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__3548\,
            I => \LED_Blink_Inst.un1_r_count_2hz_13\
        );

    \I__648\ : CascadeMux
    port map (
            O => \N__3545\,
            I => \LED_Blink_Inst.un1_r_count_2hz_20_cascade_\
        );

    \I__647\ : InMux
    port map (
            O => \N__3542\,
            I => \N__3539\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__3539\,
            I => \LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_7\
        );

    \I__645\ : InMux
    port map (
            O => \N__3536\,
            I => \N__3533\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__3533\,
            I => \LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_17\
        );

    \I__643\ : InMux
    port map (
            O => \N__3530\,
            I => \N__3524\
        );

    \I__642\ : InMux
    port map (
            O => \N__3529\,
            I => \N__3524\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__3524\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_17\
        );

    \I__640\ : InMux
    port map (
            O => \N__3521\,
            I => \LED_Blink_Inst.un6_r_count_10hz_cry_13\
        );

    \I__639\ : InMux
    port map (
            O => \N__3518\,
            I => \LED_Blink_Inst.un6_r_count_10hz_cry_14\
        );

    \I__638\ : InMux
    port map (
            O => \N__3515\,
            I => \LED_Blink_Inst.un6_r_count_10hz_cry_15\
        );

    \I__637\ : InMux
    port map (
            O => \N__3512\,
            I => \bfn_11_5_0_\
        );

    \I__636\ : InMux
    port map (
            O => \N__3509\,
            I => \LED_Blink_Inst.un6_r_count_10hz_cry_17\
        );

    \I__635\ : InMux
    port map (
            O => \N__3506\,
            I => \LED_Blink_Inst.un6_r_count_10hz_cry_18\
        );

    \I__634\ : InMux
    port map (
            O => \N__3503\,
            I => \LED_Blink_Inst.un6_r_count_10hz_cry_19\
        );

    \I__633\ : CascadeMux
    port map (
            O => \N__3500\,
            I => \LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_20_cascade_\
        );

    \I__632\ : InMux
    port map (
            O => \N__3497\,
            I => \N__3491\
        );

    \I__631\ : InMux
    port map (
            O => \N__3496\,
            I => \N__3491\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__3491\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_20\
        );

    \I__629\ : CascadeMux
    port map (
            O => \N__3488\,
            I => \N__3485\
        );

    \I__628\ : InMux
    port map (
            O => \N__3485\,
            I => \N__3479\
        );

    \I__627\ : InMux
    port map (
            O => \N__3484\,
            I => \N__3479\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__3479\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_19\
        );

    \I__625\ : InMux
    port map (
            O => \N__3476\,
            I => \N__3470\
        );

    \I__624\ : InMux
    port map (
            O => \N__3475\,
            I => \N__3470\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__3470\,
            I => \LED_Blink_Inst.r_Count_10HZZ0Z_18\
        );

    \I__622\ : InMux
    port map (
            O => \N__3467\,
            I => \LED_Blink_Inst.un6_r_count_10hz_cry_4\
        );

    \I__621\ : InMux
    port map (
            O => \N__3464\,
            I => \LED_Blink_Inst.un6_r_count_10hz_cry_5\
        );

    \I__620\ : InMux
    port map (
            O => \N__3461\,
            I => \LED_Blink_Inst.un6_r_count_10hz_cry_6\
        );

    \I__619\ : InMux
    port map (
            O => \N__3458\,
            I => \LED_Blink_Inst.un6_r_count_10hz_cry_7\
        );

    \I__618\ : InMux
    port map (
            O => \N__3455\,
            I => \bfn_11_4_0_\
        );

    \I__617\ : InMux
    port map (
            O => \N__3452\,
            I => \LED_Blink_Inst.un6_r_count_10hz_cry_9\
        );

    \I__616\ : InMux
    port map (
            O => \N__3449\,
            I => \LED_Blink_Inst.un6_r_count_10hz_cry_10\
        );

    \I__615\ : InMux
    port map (
            O => \N__3446\,
            I => \LED_Blink_Inst.un6_r_count_10hz_cry_11\
        );

    \I__614\ : InMux
    port map (
            O => \N__3443\,
            I => \LED_Blink_Inst.un6_r_count_10hz_cry_12\
        );

    \I__613\ : InMux
    port map (
            O => \N__3440\,
            I => \N__3437\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__3437\,
            I => \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_18\
        );

    \I__611\ : InMux
    port map (
            O => \N__3434\,
            I => \N__3431\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__3431\,
            I => \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_21\
        );

    \I__609\ : InMux
    port map (
            O => \N__3428\,
            I => \N__3415\
        );

    \I__608\ : InMux
    port map (
            O => \N__3427\,
            I => \N__3406\
        );

    \I__607\ : InMux
    port map (
            O => \N__3426\,
            I => \N__3406\
        );

    \I__606\ : InMux
    port map (
            O => \N__3425\,
            I => \N__3406\
        );

    \I__605\ : InMux
    port map (
            O => \N__3424\,
            I => \N__3406\
        );

    \I__604\ : InMux
    port map (
            O => \N__3423\,
            I => \N__3397\
        );

    \I__603\ : InMux
    port map (
            O => \N__3422\,
            I => \N__3397\
        );

    \I__602\ : InMux
    port map (
            O => \N__3421\,
            I => \N__3397\
        );

    \I__601\ : InMux
    port map (
            O => \N__3420\,
            I => \N__3397\
        );

    \I__600\ : InMux
    port map (
            O => \N__3419\,
            I => \N__3392\
        );

    \I__599\ : InMux
    port map (
            O => \N__3418\,
            I => \N__3392\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__3415\,
            I => \LED_Blink_Inst.un1_r_count_1hz_21\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__3406\,
            I => \LED_Blink_Inst.un1_r_count_1hz_21\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__3397\,
            I => \LED_Blink_Inst.un1_r_count_1hz_21\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__3392\,
            I => \LED_Blink_Inst.un1_r_count_1hz_21\
        );

    \I__594\ : InMux
    port map (
            O => \N__3383\,
            I => \N__3380\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__3380\,
            I => \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_17\
        );

    \I__592\ : CascadeMux
    port map (
            O => \N__3377\,
            I => \N__3366\
        );

    \I__591\ : CascadeMux
    port map (
            O => \N__3376\,
            I => \N__3363\
        );

    \I__590\ : CascadeMux
    port map (
            O => \N__3375\,
            I => \N__3360\
        );

    \I__589\ : CascadeMux
    port map (
            O => \N__3374\,
            I => \N__3357\
        );

    \I__588\ : CascadeMux
    port map (
            O => \N__3373\,
            I => \N__3354\
        );

    \I__587\ : CascadeMux
    port map (
            O => \N__3372\,
            I => \N__3351\
        );

    \I__586\ : InMux
    port map (
            O => \N__3371\,
            I => \N__3347\
        );

    \I__585\ : CascadeMux
    port map (
            O => \N__3370\,
            I => \N__3342\
        );

    \I__584\ : InMux
    port map (
            O => \N__3369\,
            I => \N__3339\
        );

    \I__583\ : InMux
    port map (
            O => \N__3366\,
            I => \N__3334\
        );

    \I__582\ : InMux
    port map (
            O => \N__3363\,
            I => \N__3334\
        );

    \I__581\ : InMux
    port map (
            O => \N__3360\,
            I => \N__3329\
        );

    \I__580\ : InMux
    port map (
            O => \N__3357\,
            I => \N__3329\
        );

    \I__579\ : InMux
    port map (
            O => \N__3354\,
            I => \N__3326\
        );

    \I__578\ : InMux
    port map (
            O => \N__3351\,
            I => \N__3321\
        );

    \I__577\ : InMux
    port map (
            O => \N__3350\,
            I => \N__3321\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__3347\,
            I => \N__3318\
        );

    \I__575\ : InMux
    port map (
            O => \N__3346\,
            I => \N__3311\
        );

    \I__574\ : InMux
    port map (
            O => \N__3345\,
            I => \N__3311\
        );

    \I__573\ : InMux
    port map (
            O => \N__3342\,
            I => \N__3311\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__3339\,
            I => \N__3308\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__3334\,
            I => \N__3303\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__3329\,
            I => \N__3303\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__3326\,
            I => \N__3296\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__3321\,
            I => \N__3296\
        );

    \I__567\ : Span4Mux_h
    port map (
            O => \N__3318\,
            I => \N__3296\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__3311\,
            I => \LED_Blink_Inst.un1_r_count_1hz_17\
        );

    \I__565\ : Odrv4
    port map (
            O => \N__3308\,
            I => \LED_Blink_Inst.un1_r_count_1hz_17\
        );

    \I__564\ : Odrv12
    port map (
            O => \N__3303\,
            I => \LED_Blink_Inst.un1_r_count_1hz_17\
        );

    \I__563\ : Odrv4
    port map (
            O => \N__3296\,
            I => \LED_Blink_Inst.un1_r_count_1hz_17\
        );

    \I__562\ : InMux
    port map (
            O => \N__3287\,
            I => \N__3270\
        );

    \I__561\ : InMux
    port map (
            O => \N__3286\,
            I => \N__3270\
        );

    \I__560\ : InMux
    port map (
            O => \N__3285\,
            I => \N__3270\
        );

    \I__559\ : InMux
    port map (
            O => \N__3284\,
            I => \N__3270\
        );

    \I__558\ : InMux
    port map (
            O => \N__3283\,
            I => \N__3265\
        );

    \I__557\ : InMux
    port map (
            O => \N__3282\,
            I => \N__3256\
        );

    \I__556\ : InMux
    port map (
            O => \N__3281\,
            I => \N__3256\
        );

    \I__555\ : InMux
    port map (
            O => \N__3280\,
            I => \N__3256\
        );

    \I__554\ : InMux
    port map (
            O => \N__3279\,
            I => \N__3256\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__3270\,
            I => \N__3253\
        );

    \I__552\ : InMux
    port map (
            O => \N__3269\,
            I => \N__3248\
        );

    \I__551\ : InMux
    port map (
            O => \N__3268\,
            I => \N__3248\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__3265\,
            I => \LED_Blink_Inst.un1_r_count_1hz_16\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__3256\,
            I => \LED_Blink_Inst.un1_r_count_1hz_16\
        );

    \I__548\ : Odrv4
    port map (
            O => \N__3253\,
            I => \LED_Blink_Inst.un1_r_count_1hz_16\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__3248\,
            I => \LED_Blink_Inst.un1_r_count_1hz_16\
        );

    \I__546\ : InMux
    port map (
            O => \N__3239\,
            I => \N__3235\
        );

    \I__545\ : InMux
    port map (
            O => \N__3238\,
            I => \N__3232\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__3235\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_20\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__3232\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_20\
        );

    \I__542\ : InMux
    port map (
            O => \N__3227\,
            I => \N__3223\
        );

    \I__541\ : InMux
    port map (
            O => \N__3226\,
            I => \N__3220\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__3223\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_18\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__3220\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_18\
        );

    \I__538\ : CascadeMux
    port map (
            O => \N__3215\,
            I => \N__3211\
        );

    \I__537\ : InMux
    port map (
            O => \N__3214\,
            I => \N__3208\
        );

    \I__536\ : InMux
    port map (
            O => \N__3211\,
            I => \N__3205\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__3208\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_21\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__3205\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_21\
        );

    \I__533\ : InMux
    port map (
            O => \N__3200\,
            I => \N__3196\
        );

    \I__532\ : InMux
    port map (
            O => \N__3199\,
            I => \N__3193\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__3196\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_17\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__3193\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_17\
        );

    \I__529\ : InMux
    port map (
            O => \N__3188\,
            I => \N__3185\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__3185\,
            I => \LED_Blink_Inst.un1_r_count_1hz_15\
        );

    \I__527\ : InMux
    port map (
            O => \N__3182\,
            I => \LED_Blink_Inst.un6_r_count_10hz_cry_1\
        );

    \I__526\ : InMux
    port map (
            O => \N__3179\,
            I => \LED_Blink_Inst.un6_r_count_10hz_cry_2\
        );

    \I__525\ : InMux
    port map (
            O => \N__3176\,
            I => \LED_Blink_Inst.un6_r_count_10hz_cry_3\
        );

    \I__524\ : InMux
    port map (
            O => \N__3173\,
            I => \N__3166\
        );

    \I__523\ : InMux
    port map (
            O => \N__3172\,
            I => \N__3166\
        );

    \I__522\ : InMux
    port map (
            O => \N__3171\,
            I => \N__3163\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__3166\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_1\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__3163\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_1\
        );

    \I__519\ : CascadeMux
    port map (
            O => \N__3158\,
            I => \N__3155\
        );

    \I__518\ : InMux
    port map (
            O => \N__3155\,
            I => \N__3152\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__3152\,
            I => \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_11\
        );

    \I__516\ : InMux
    port map (
            O => \N__3149\,
            I => \N__3145\
        );

    \I__515\ : InMux
    port map (
            O => \N__3148\,
            I => \N__3142\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__3145\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_11\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__3142\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_11\
        );

    \I__512\ : InMux
    port map (
            O => \N__3137\,
            I => \N__3134\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__3134\,
            I => \N__3131\
        );

    \I__510\ : Odrv4
    port map (
            O => \N__3131\,
            I => \LED_Blink_Inst.un1_r_count_1hz_13\
        );

    \I__509\ : CascadeMux
    port map (
            O => \N__3128\,
            I => \LED_Blink_Inst.un1_r_count_1hz_14_cascade_\
        );

    \I__508\ : InMux
    port map (
            O => \N__3125\,
            I => \N__3122\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__3122\,
            I => \LED_Blink_Inst.un1_r_count_1hz_12\
        );

    \I__506\ : CascadeMux
    port map (
            O => \N__3119\,
            I => \LED_Blink_Inst.un1_r_count_1hz_21_cascade_\
        );

    \I__505\ : InMux
    port map (
            O => \N__3116\,
            I => \N__3113\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__3113\,
            I => \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_12\
        );

    \I__503\ : InMux
    port map (
            O => \N__3110\,
            I => \N__3106\
        );

    \I__502\ : InMux
    port map (
            O => \N__3109\,
            I => \N__3103\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__3106\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_12\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__3103\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_12\
        );

    \I__499\ : InMux
    port map (
            O => \N__3098\,
            I => \N__3094\
        );

    \I__498\ : InMux
    port map (
            O => \N__3097\,
            I => \N__3091\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__3094\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_22\
        );

    \I__496\ : LocalMux
    port map (
            O => \N__3091\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_22\
        );

    \I__495\ : InMux
    port map (
            O => \N__3086\,
            I => \N__3082\
        );

    \I__494\ : InMux
    port map (
            O => \N__3085\,
            I => \N__3079\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__3082\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_19\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__3079\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_19\
        );

    \I__491\ : CascadeMux
    port map (
            O => \N__3074\,
            I => \N__3071\
        );

    \I__490\ : InMux
    port map (
            O => \N__3071\,
            I => \N__3067\
        );

    \I__489\ : InMux
    port map (
            O => \N__3070\,
            I => \N__3064\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__3067\,
            I => \N__3061\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__3064\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_23\
        );

    \I__486\ : Odrv4
    port map (
            O => \N__3061\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_23\
        );

    \I__485\ : InMux
    port map (
            O => \N__3056\,
            I => \N__3052\
        );

    \I__484\ : InMux
    port map (
            O => \N__3055\,
            I => \N__3049\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__3052\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_14\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__3049\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_14\
        );

    \I__481\ : CascadeMux
    port map (
            O => \N__3044\,
            I => \LED_Blink_Inst.un1_r_count_1hz_16_cascade_\
        );

    \I__480\ : InMux
    port map (
            O => \N__3041\,
            I => \N__3038\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__3038\,
            I => \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_16\
        );

    \I__478\ : CascadeMux
    port map (
            O => \N__3035\,
            I => \N__3032\
        );

    \I__477\ : InMux
    port map (
            O => \N__3032\,
            I => \N__3028\
        );

    \I__476\ : InMux
    port map (
            O => \N__3031\,
            I => \N__3025\
        );

    \I__475\ : LocalMux
    port map (
            O => \N__3028\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_16\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__3025\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_16\
        );

    \I__473\ : InMux
    port map (
            O => \N__3020\,
            I => \N__3017\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__3017\,
            I => \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_9\
        );

    \I__471\ : InMux
    port map (
            O => \N__3014\,
            I => \N__3010\
        );

    \I__470\ : InMux
    port map (
            O => \N__3013\,
            I => \N__3007\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__3010\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_9\
        );

    \I__468\ : LocalMux
    port map (
            O => \N__3007\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_9\
        );

    \I__467\ : InMux
    port map (
            O => \N__3002\,
            I => \N__2999\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__2999\,
            I => \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_20\
        );

    \I__465\ : InMux
    port map (
            O => \N__2996\,
            I => \LED_Blink_Inst.un4_r_count_1hz_cry_22\
        );

    \I__464\ : CascadeMux
    port map (
            O => \N__2993\,
            I => \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_23_cascade_\
        );

    \I__463\ : InMux
    port map (
            O => \N__2990\,
            I => \N__2987\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__2987\,
            I => \N__2983\
        );

    \I__461\ : InMux
    port map (
            O => \N__2986\,
            I => \N__2980\
        );

    \I__460\ : Odrv4
    port map (
            O => \N__2983\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_13\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__2980\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_13\
        );

    \I__458\ : InMux
    port map (
            O => \N__2975\,
            I => \N__2972\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__2972\,
            I => \N__2968\
        );

    \I__456\ : InMux
    port map (
            O => \N__2971\,
            I => \N__2965\
        );

    \I__455\ : Odrv4
    port map (
            O => \N__2968\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_10\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__2965\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_10\
        );

    \I__453\ : CascadeMux
    port map (
            O => \N__2960\,
            I => \N__2957\
        );

    \I__452\ : InMux
    port map (
            O => \N__2957\,
            I => \N__2953\
        );

    \I__451\ : CascadeMux
    port map (
            O => \N__2956\,
            I => \N__2950\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__2953\,
            I => \N__2947\
        );

    \I__449\ : InMux
    port map (
            O => \N__2950\,
            I => \N__2944\
        );

    \I__448\ : Odrv4
    port map (
            O => \N__2947\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_15\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__2944\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_15\
        );

    \I__446\ : InMux
    port map (
            O => \N__2939\,
            I => \N__2936\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__2936\,
            I => \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_8\
        );

    \I__444\ : IoInMux
    port map (
            O => \N__2933\,
            I => \N__2930\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__2930\,
            I => \N__2926\
        );

    \I__442\ : CascadeMux
    port map (
            O => \N__2929\,
            I => \N__2923\
        );

    \I__441\ : Span4Mux_s2_h
    port map (
            O => \N__2926\,
            I => \N__2920\
        );

    \I__440\ : InMux
    port map (
            O => \N__2923\,
            I => \N__2917\
        );

    \I__439\ : Odrv4
    port map (
            O => \N__2920\,
            I => \o_LED_4_c\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__2917\,
            I => \o_LED_4_c\
        );

    \I__437\ : InMux
    port map (
            O => \N__2912\,
            I => \N__2908\
        );

    \I__436\ : InMux
    port map (
            O => \N__2911\,
            I => \N__2905\
        );

    \I__435\ : LocalMux
    port map (
            O => \N__2908\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_5\
        );

    \I__434\ : LocalMux
    port map (
            O => \N__2905\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_5\
        );

    \I__433\ : InMux
    port map (
            O => \N__2900\,
            I => \N__2896\
        );

    \I__432\ : InMux
    port map (
            O => \N__2899\,
            I => \N__2893\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__2896\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_6\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__2893\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_6\
        );

    \I__429\ : CascadeMux
    port map (
            O => \N__2888\,
            I => \N__2885\
        );

    \I__428\ : InMux
    port map (
            O => \N__2885\,
            I => \N__2881\
        );

    \I__427\ : InMux
    port map (
            O => \N__2884\,
            I => \N__2878\
        );

    \I__426\ : LocalMux
    port map (
            O => \N__2881\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_7\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__2878\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_7\
        );

    \I__424\ : InMux
    port map (
            O => \N__2873\,
            I => \N__2869\
        );

    \I__423\ : InMux
    port map (
            O => \N__2872\,
            I => \N__2866\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__2869\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_4\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__2866\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_4\
        );

    \I__420\ : CascadeMux
    port map (
            O => \N__2861\,
            I => \N__2857\
        );

    \I__419\ : CascadeMux
    port map (
            O => \N__2860\,
            I => \N__2852\
        );

    \I__418\ : InMux
    port map (
            O => \N__2857\,
            I => \N__2847\
        );

    \I__417\ : InMux
    port map (
            O => \N__2856\,
            I => \N__2847\
        );

    \I__416\ : InMux
    port map (
            O => \N__2855\,
            I => \N__2844\
        );

    \I__415\ : InMux
    port map (
            O => \N__2852\,
            I => \N__2841\
        );

    \I__414\ : LocalMux
    port map (
            O => \N__2847\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_0\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__2844\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_0\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__2841\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_0\
        );

    \I__411\ : InMux
    port map (
            O => \N__2834\,
            I => \N__2830\
        );

    \I__410\ : InMux
    port map (
            O => \N__2833\,
            I => \N__2827\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__2830\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_3\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__2827\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_3\
        );

    \I__407\ : InMux
    port map (
            O => \N__2822\,
            I => \N__2818\
        );

    \I__406\ : InMux
    port map (
            O => \N__2821\,
            I => \N__2815\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__2818\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_2\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__2815\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_2\
        );

    \I__403\ : CascadeMux
    port map (
            O => \N__2810\,
            I => \N__2807\
        );

    \I__402\ : InMux
    port map (
            O => \N__2807\,
            I => \N__2803\
        );

    \I__401\ : InMux
    port map (
            O => \N__2806\,
            I => \N__2800\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__2803\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_8\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__2800\,
            I => \LED_Blink_Inst.r_Count_1HZZ0Z_8\
        );

    \I__398\ : InMux
    port map (
            O => \N__2795\,
            I => \LED_Blink_Inst.un4_r_count_1hz_cry_13\
        );

    \I__397\ : InMux
    port map (
            O => \N__2792\,
            I => \LED_Blink_Inst.un4_r_count_1hz_cry_14\
        );

    \I__396\ : InMux
    port map (
            O => \N__2789\,
            I => \LED_Blink_Inst.un4_r_count_1hz_cry_15\
        );

    \I__395\ : InMux
    port map (
            O => \N__2786\,
            I => \bfn_8_9_0_\
        );

    \I__394\ : InMux
    port map (
            O => \N__2783\,
            I => \LED_Blink_Inst.un4_r_count_1hz_cry_17\
        );

    \I__393\ : InMux
    port map (
            O => \N__2780\,
            I => \LED_Blink_Inst.un4_r_count_1hz_cry_18\
        );

    \I__392\ : InMux
    port map (
            O => \N__2777\,
            I => \LED_Blink_Inst.un4_r_count_1hz_cry_19\
        );

    \I__391\ : InMux
    port map (
            O => \N__2774\,
            I => \LED_Blink_Inst.un4_r_count_1hz_cry_20\
        );

    \I__390\ : InMux
    port map (
            O => \N__2771\,
            I => \LED_Blink_Inst.un4_r_count_1hz_cry_21\
        );

    \I__389\ : InMux
    port map (
            O => \N__2768\,
            I => \LED_Blink_Inst.un4_r_count_1hz_cry_4\
        );

    \I__388\ : InMux
    port map (
            O => \N__2765\,
            I => \LED_Blink_Inst.un4_r_count_1hz_cry_5\
        );

    \I__387\ : InMux
    port map (
            O => \N__2762\,
            I => \LED_Blink_Inst.un4_r_count_1hz_cry_6\
        );

    \I__386\ : InMux
    port map (
            O => \N__2759\,
            I => \LED_Blink_Inst.un4_r_count_1hz_cry_7\
        );

    \I__385\ : InMux
    port map (
            O => \N__2756\,
            I => \bfn_8_8_0_\
        );

    \I__384\ : InMux
    port map (
            O => \N__2753\,
            I => \LED_Blink_Inst.un4_r_count_1hz_cry_9\
        );

    \I__383\ : InMux
    port map (
            O => \N__2750\,
            I => \LED_Blink_Inst.un4_r_count_1hz_cry_10\
        );

    \I__382\ : InMux
    port map (
            O => \N__2747\,
            I => \LED_Blink_Inst.un4_r_count_1hz_cry_11\
        );

    \I__381\ : InMux
    port map (
            O => \N__2744\,
            I => \LED_Blink_Inst.un4_r_count_1hz_cry_12\
        );

    \I__380\ : InMux
    port map (
            O => \N__2741\,
            I => \N__2738\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__2738\,
            I => \LED_Blink_Inst.un1_r_count_5hz_11\
        );

    \I__378\ : InMux
    port map (
            O => \N__2735\,
            I => \N__2731\
        );

    \I__377\ : InMux
    port map (
            O => \N__2734\,
            I => \N__2728\
        );

    \I__376\ : LocalMux
    port map (
            O => \N__2731\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_11\
        );

    \I__375\ : LocalMux
    port map (
            O => \N__2728\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_11\
        );

    \I__374\ : CascadeMux
    port map (
            O => \N__2723\,
            I => \LED_Blink_Inst.un1_r_count_5hz_17_cascade_\
        );

    \I__373\ : CascadeMux
    port map (
            O => \N__2720\,
            I => \N__2714\
        );

    \I__372\ : InMux
    port map (
            O => \N__2719\,
            I => \N__2711\
        );

    \I__371\ : InMux
    port map (
            O => \N__2718\,
            I => \N__2706\
        );

    \I__370\ : InMux
    port map (
            O => \N__2717\,
            I => \N__2706\
        );

    \I__369\ : InMux
    port map (
            O => \N__2714\,
            I => \N__2703\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__2711\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_0\
        );

    \I__367\ : LocalMux
    port map (
            O => \N__2706\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_0\
        );

    \I__366\ : LocalMux
    port map (
            O => \N__2703\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_0\
        );

    \I__365\ : CascadeMux
    port map (
            O => \N__2696\,
            I => \LED_Blink_Inst.un1_r_count_5hz_19_cascade_\
        );

    \I__364\ : InMux
    port map (
            O => \N__2693\,
            I => \N__2690\
        );

    \I__363\ : LocalMux
    port map (
            O => \N__2690\,
            I => \LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_17\
        );

    \I__362\ : CascadeMux
    port map (
            O => \N__2687\,
            I => \N__2684\
        );

    \I__361\ : InMux
    port map (
            O => \N__2684\,
            I => \N__2680\
        );

    \I__360\ : InMux
    port map (
            O => \N__2683\,
            I => \N__2677\
        );

    \I__359\ : LocalMux
    port map (
            O => \N__2680\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_17\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__2677\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_17\
        );

    \I__357\ : InMux
    port map (
            O => \N__2672\,
            I => \N__2668\
        );

    \I__356\ : InMux
    port map (
            O => \N__2671\,
            I => \N__2665\
        );

    \I__355\ : LocalMux
    port map (
            O => \N__2668\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_9\
        );

    \I__354\ : LocalMux
    port map (
            O => \N__2665\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_9\
        );

    \I__353\ : InMux
    port map (
            O => \N__2660\,
            I => \N__2656\
        );

    \I__352\ : InMux
    port map (
            O => \N__2659\,
            I => \N__2653\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__2656\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_14\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__2653\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_14\
        );

    \I__349\ : CascadeMux
    port map (
            O => \N__2648\,
            I => \N__2645\
        );

    \I__348\ : InMux
    port map (
            O => \N__2645\,
            I => \N__2641\
        );

    \I__347\ : InMux
    port map (
            O => \N__2644\,
            I => \N__2638\
        );

    \I__346\ : LocalMux
    port map (
            O => \N__2641\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_16\
        );

    \I__345\ : LocalMux
    port map (
            O => \N__2638\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_16\
        );

    \I__344\ : InMux
    port map (
            O => \N__2633\,
            I => \N__2629\
        );

    \I__343\ : InMux
    port map (
            O => \N__2632\,
            I => \N__2626\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__2629\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_12\
        );

    \I__341\ : LocalMux
    port map (
            O => \N__2626\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_12\
        );

    \I__340\ : CascadeMux
    port map (
            O => \N__2621\,
            I => \N__2613\
        );

    \I__339\ : InMux
    port map (
            O => \N__2620\,
            I => \N__2609\
        );

    \I__338\ : CascadeMux
    port map (
            O => \N__2619\,
            I => \N__2606\
        );

    \I__337\ : InMux
    port map (
            O => \N__2618\,
            I => \N__2597\
        );

    \I__336\ : InMux
    port map (
            O => \N__2617\,
            I => \N__2597\
        );

    \I__335\ : InMux
    port map (
            O => \N__2616\,
            I => \N__2597\
        );

    \I__334\ : InMux
    port map (
            O => \N__2613\,
            I => \N__2597\
        );

    \I__333\ : CascadeMux
    port map (
            O => \N__2612\,
            I => \N__2592\
        );

    \I__332\ : LocalMux
    port map (
            O => \N__2609\,
            I => \N__2589\
        );

    \I__331\ : InMux
    port map (
            O => \N__2606\,
            I => \N__2586\
        );

    \I__330\ : LocalMux
    port map (
            O => \N__2597\,
            I => \N__2583\
        );

    \I__329\ : InMux
    port map (
            O => \N__2596\,
            I => \N__2578\
        );

    \I__328\ : InMux
    port map (
            O => \N__2595\,
            I => \N__2578\
        );

    \I__327\ : InMux
    port map (
            O => \N__2592\,
            I => \N__2575\
        );

    \I__326\ : Odrv4
    port map (
            O => \N__2589\,
            I => \LED_Blink_Inst.un1_r_count_5hz_15\
        );

    \I__325\ : LocalMux
    port map (
            O => \N__2586\,
            I => \LED_Blink_Inst.un1_r_count_5hz_15\
        );

    \I__324\ : Odrv4
    port map (
            O => \N__2583\,
            I => \LED_Blink_Inst.un1_r_count_5hz_15\
        );

    \I__323\ : LocalMux
    port map (
            O => \N__2578\,
            I => \LED_Blink_Inst.un1_r_count_5hz_15\
        );

    \I__322\ : LocalMux
    port map (
            O => \N__2575\,
            I => \LED_Blink_Inst.un1_r_count_5hz_15\
        );

    \I__321\ : CascadeMux
    port map (
            O => \N__2564\,
            I => \N__2557\
        );

    \I__320\ : CascadeMux
    port map (
            O => \N__2563\,
            I => \N__2552\
        );

    \I__319\ : CascadeMux
    port map (
            O => \N__2562\,
            I => \N__2549\
        );

    \I__318\ : CascadeMux
    port map (
            O => \N__2561\,
            I => \N__2545\
        );

    \I__317\ : InMux
    port map (
            O => \N__2560\,
            I => \N__2539\
        );

    \I__316\ : InMux
    port map (
            O => \N__2557\,
            I => \N__2539\
        );

    \I__315\ : InMux
    port map (
            O => \N__2556\,
            I => \N__2530\
        );

    \I__314\ : InMux
    port map (
            O => \N__2555\,
            I => \N__2530\
        );

    \I__313\ : InMux
    port map (
            O => \N__2552\,
            I => \N__2530\
        );

    \I__312\ : InMux
    port map (
            O => \N__2549\,
            I => \N__2530\
        );

    \I__311\ : InMux
    port map (
            O => \N__2548\,
            I => \N__2523\
        );

    \I__310\ : InMux
    port map (
            O => \N__2545\,
            I => \N__2523\
        );

    \I__309\ : InMux
    port map (
            O => \N__2544\,
            I => \N__2523\
        );

    \I__308\ : LocalMux
    port map (
            O => \N__2539\,
            I => \LED_Blink_Inst.un1_r_count_5hz_19\
        );

    \I__307\ : LocalMux
    port map (
            O => \N__2530\,
            I => \LED_Blink_Inst.un1_r_count_5hz_19\
        );

    \I__306\ : LocalMux
    port map (
            O => \N__2523\,
            I => \LED_Blink_Inst.un1_r_count_5hz_19\
        );

    \I__305\ : InMux
    port map (
            O => \N__2516\,
            I => \N__2504\
        );

    \I__304\ : InMux
    port map (
            O => \N__2515\,
            I => \N__2504\
        );

    \I__303\ : InMux
    port map (
            O => \N__2514\,
            I => \N__2504\
        );

    \I__302\ : InMux
    port map (
            O => \N__2513\,
            I => \N__2504\
        );

    \I__301\ : LocalMux
    port map (
            O => \N__2504\,
            I => \N__2495\
        );

    \I__300\ : InMux
    port map (
            O => \N__2503\,
            I => \N__2486\
        );

    \I__299\ : InMux
    port map (
            O => \N__2502\,
            I => \N__2486\
        );

    \I__298\ : InMux
    port map (
            O => \N__2501\,
            I => \N__2486\
        );

    \I__297\ : InMux
    port map (
            O => \N__2500\,
            I => \N__2486\
        );

    \I__296\ : InMux
    port map (
            O => \N__2499\,
            I => \N__2481\
        );

    \I__295\ : InMux
    port map (
            O => \N__2498\,
            I => \N__2481\
        );

    \I__294\ : Odrv4
    port map (
            O => \N__2495\,
            I => \LED_Blink_Inst.un1_r_count_5hz_14\
        );

    \I__293\ : LocalMux
    port map (
            O => \N__2486\,
            I => \LED_Blink_Inst.un1_r_count_5hz_14\
        );

    \I__292\ : LocalMux
    port map (
            O => \N__2481\,
            I => \LED_Blink_Inst.un1_r_count_5hz_14\
        );

    \I__291\ : CascadeMux
    port map (
            O => \N__2474\,
            I => \LED_Blink_Inst.un1_r_count_5hz_15_cascade_\
        );

    \I__290\ : InMux
    port map (
            O => \N__2471\,
            I => \N__2468\
        );

    \I__289\ : LocalMux
    port map (
            O => \N__2468\,
            I => \LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_10\
        );

    \I__288\ : InMux
    port map (
            O => \N__2465\,
            I => \N__2461\
        );

    \I__287\ : InMux
    port map (
            O => \N__2464\,
            I => \N__2458\
        );

    \I__286\ : LocalMux
    port map (
            O => \N__2461\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_10\
        );

    \I__285\ : LocalMux
    port map (
            O => \N__2458\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_10\
        );

    \I__284\ : InMux
    port map (
            O => \N__2453\,
            I => \LED_Blink_Inst.un4_r_count_1hz_cry_1\
        );

    \I__283\ : InMux
    port map (
            O => \N__2450\,
            I => \LED_Blink_Inst.un4_r_count_1hz_cry_2\
        );

    \I__282\ : InMux
    port map (
            O => \N__2447\,
            I => \LED_Blink_Inst.un4_r_count_1hz_cry_3\
        );

    \I__281\ : InMux
    port map (
            O => \N__2444\,
            I => \N__2440\
        );

    \I__280\ : InMux
    port map (
            O => \N__2443\,
            I => \N__2437\
        );

    \I__279\ : LocalMux
    port map (
            O => \N__2440\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_4\
        );

    \I__278\ : LocalMux
    port map (
            O => \N__2437\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_4\
        );

    \I__277\ : InMux
    port map (
            O => \N__2432\,
            I => \N__2428\
        );

    \I__276\ : InMux
    port map (
            O => \N__2431\,
            I => \N__2425\
        );

    \I__275\ : LocalMux
    port map (
            O => \N__2428\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_2\
        );

    \I__274\ : LocalMux
    port map (
            O => \N__2425\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_2\
        );

    \I__273\ : CascadeMux
    port map (
            O => \N__2420\,
            I => \N__2417\
        );

    \I__272\ : InMux
    port map (
            O => \N__2417\,
            I => \N__2413\
        );

    \I__271\ : InMux
    port map (
            O => \N__2416\,
            I => \N__2410\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__2413\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_6\
        );

    \I__269\ : LocalMux
    port map (
            O => \N__2410\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_6\
        );

    \I__268\ : InMux
    port map (
            O => \N__2405\,
            I => \N__2401\
        );

    \I__267\ : InMux
    port map (
            O => \N__2404\,
            I => \N__2398\
        );

    \I__266\ : LocalMux
    port map (
            O => \N__2401\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_7\
        );

    \I__265\ : LocalMux
    port map (
            O => \N__2398\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_7\
        );

    \I__264\ : InMux
    port map (
            O => \N__2393\,
            I => \N__2386\
        );

    \I__263\ : InMux
    port map (
            O => \N__2392\,
            I => \N__2386\
        );

    \I__262\ : InMux
    port map (
            O => \N__2391\,
            I => \N__2383\
        );

    \I__261\ : LocalMux
    port map (
            O => \N__2386\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_1\
        );

    \I__260\ : LocalMux
    port map (
            O => \N__2383\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_1\
        );

    \I__259\ : InMux
    port map (
            O => \N__2378\,
            I => \N__2375\
        );

    \I__258\ : LocalMux
    port map (
            O => \N__2375\,
            I => \LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_8\
        );

    \I__257\ : InMux
    port map (
            O => \N__2372\,
            I => \N__2368\
        );

    \I__256\ : InMux
    port map (
            O => \N__2371\,
            I => \N__2365\
        );

    \I__255\ : LocalMux
    port map (
            O => \N__2368\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_8\
        );

    \I__254\ : LocalMux
    port map (
            O => \N__2365\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_8\
        );

    \I__253\ : IoInMux
    port map (
            O => \N__2360\,
            I => \N__2357\
        );

    \I__252\ : LocalMux
    port map (
            O => \N__2357\,
            I => \N__2353\
        );

    \I__251\ : CascadeMux
    port map (
            O => \N__2356\,
            I => \N__2350\
        );

    \I__250\ : Span4Mux_s3_h
    port map (
            O => \N__2353\,
            I => \N__2347\
        );

    \I__249\ : InMux
    port map (
            O => \N__2350\,
            I => \N__2344\
        );

    \I__248\ : Odrv4
    port map (
            O => \N__2347\,
            I => \o_LED_2_c\
        );

    \I__247\ : LocalMux
    port map (
            O => \N__2344\,
            I => \o_LED_2_c\
        );

    \I__246\ : InMux
    port map (
            O => \N__2339\,
            I => \N__2336\
        );

    \I__245\ : LocalMux
    port map (
            O => \N__2336\,
            I => \LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_13\
        );

    \I__244\ : InMux
    port map (
            O => \N__2333\,
            I => \N__2329\
        );

    \I__243\ : InMux
    port map (
            O => \N__2332\,
            I => \N__2326\
        );

    \I__242\ : LocalMux
    port map (
            O => \N__2329\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_13\
        );

    \I__241\ : LocalMux
    port map (
            O => \N__2326\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_13\
        );

    \I__240\ : InMux
    port map (
            O => \N__2321\,
            I => \N__2317\
        );

    \I__239\ : InMux
    port map (
            O => \N__2320\,
            I => \N__2314\
        );

    \I__238\ : LocalMux
    port map (
            O => \N__2317\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_18\
        );

    \I__237\ : LocalMux
    port map (
            O => \N__2314\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_18\
        );

    \I__236\ : InMux
    port map (
            O => \N__2309\,
            I => \N__2305\
        );

    \I__235\ : InMux
    port map (
            O => \N__2308\,
            I => \N__2302\
        );

    \I__234\ : LocalMux
    port map (
            O => \N__2305\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_5\
        );

    \I__233\ : LocalMux
    port map (
            O => \N__2302\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_5\
        );

    \I__232\ : InMux
    port map (
            O => \N__2297\,
            I => \N__2293\
        );

    \I__231\ : InMux
    port map (
            O => \N__2296\,
            I => \N__2290\
        );

    \I__230\ : LocalMux
    port map (
            O => \N__2293\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_3\
        );

    \I__229\ : LocalMux
    port map (
            O => \N__2290\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_3\
        );

    \I__228\ : CascadeMux
    port map (
            O => \N__2285\,
            I => \LED_Blink_Inst.un1_r_count_5hz_13_cascade_\
        );

    \I__227\ : InMux
    port map (
            O => \N__2282\,
            I => \N__2279\
        );

    \I__226\ : LocalMux
    port map (
            O => \N__2279\,
            I => \LED_Blink_Inst.un1_r_count_5hz_3\
        );

    \I__225\ : InMux
    port map (
            O => \N__2276\,
            I => \LED_Blink_Inst.un4_r_count_5hz_cry_17\
        );

    \I__224\ : InMux
    port map (
            O => \N__2273\,
            I => \LED_Blink_Inst.un4_r_count_5hz_cry_18\
        );

    \I__223\ : InMux
    port map (
            O => \N__2270\,
            I => \LED_Blink_Inst.un4_r_count_5hz_cry_19\
        );

    \I__222\ : InMux
    port map (
            O => \N__2267\,
            I => \LED_Blink_Inst.un4_r_count_5hz_cry_20\
        );

    \I__221\ : InMux
    port map (
            O => \N__2264\,
            I => \N__2261\
        );

    \I__220\ : LocalMux
    port map (
            O => \N__2261\,
            I => \LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_18\
        );

    \I__219\ : InMux
    port map (
            O => \N__2258\,
            I => \N__2255\
        );

    \I__218\ : LocalMux
    port map (
            O => \N__2255\,
            I => \LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_21\
        );

    \I__217\ : InMux
    port map (
            O => \N__2252\,
            I => \N__2246\
        );

    \I__216\ : InMux
    port map (
            O => \N__2251\,
            I => \N__2246\
        );

    \I__215\ : LocalMux
    port map (
            O => \N__2246\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_19\
        );

    \I__214\ : InMux
    port map (
            O => \N__2243\,
            I => \N__2237\
        );

    \I__213\ : InMux
    port map (
            O => \N__2242\,
            I => \N__2237\
        );

    \I__212\ : LocalMux
    port map (
            O => \N__2237\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_20\
        );

    \I__211\ : CascadeMux
    port map (
            O => \N__2234\,
            I => \N__2230\
        );

    \I__210\ : InMux
    port map (
            O => \N__2233\,
            I => \N__2225\
        );

    \I__209\ : InMux
    port map (
            O => \N__2230\,
            I => \N__2225\
        );

    \I__208\ : LocalMux
    port map (
            O => \N__2225\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_21\
        );

    \I__207\ : InMux
    port map (
            O => \N__2222\,
            I => \N__2218\
        );

    \I__206\ : InMux
    port map (
            O => \N__2221\,
            I => \N__2215\
        );

    \I__205\ : LocalMux
    port map (
            O => \N__2218\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_15\
        );

    \I__204\ : LocalMux
    port map (
            O => \N__2215\,
            I => \LED_Blink_Inst.r_Count_5HZZ0Z_15\
        );

    \I__203\ : InMux
    port map (
            O => \N__2210\,
            I => \N__2207\
        );

    \I__202\ : LocalMux
    port map (
            O => \N__2207\,
            I => \LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_7\
        );

    \I__201\ : InMux
    port map (
            O => \N__2204\,
            I => \N__2201\
        );

    \I__200\ : LocalMux
    port map (
            O => \N__2201\,
            I => \LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_5\
        );

    \I__199\ : InMux
    port map (
            O => \N__2198\,
            I => \bfn_7_6_0_\
        );

    \I__198\ : InMux
    port map (
            O => \N__2195\,
            I => \LED_Blink_Inst.un4_r_count_5hz_cry_9\
        );

    \I__197\ : InMux
    port map (
            O => \N__2192\,
            I => \LED_Blink_Inst.un4_r_count_5hz_cry_10\
        );

    \I__196\ : InMux
    port map (
            O => \N__2189\,
            I => \LED_Blink_Inst.un4_r_count_5hz_cry_11\
        );

    \I__195\ : InMux
    port map (
            O => \N__2186\,
            I => \LED_Blink_Inst.un4_r_count_5hz_cry_12\
        );

    \I__194\ : InMux
    port map (
            O => \N__2183\,
            I => \LED_Blink_Inst.un4_r_count_5hz_cry_13\
        );

    \I__193\ : InMux
    port map (
            O => \N__2180\,
            I => \LED_Blink_Inst.un4_r_count_5hz_cry_14\
        );

    \I__192\ : InMux
    port map (
            O => \N__2177\,
            I => \LED_Blink_Inst.un4_r_count_5hz_cry_15\
        );

    \I__191\ : InMux
    port map (
            O => \N__2174\,
            I => \bfn_7_7_0_\
        );

    \I__190\ : InMux
    port map (
            O => \N__2171\,
            I => \LED_Blink_Inst.un4_r_count_5hz_cry_1\
        );

    \I__189\ : InMux
    port map (
            O => \N__2168\,
            I => \LED_Blink_Inst.un4_r_count_5hz_cry_2\
        );

    \I__188\ : InMux
    port map (
            O => \N__2165\,
            I => \LED_Blink_Inst.un4_r_count_5hz_cry_3\
        );

    \I__187\ : InMux
    port map (
            O => \N__2162\,
            I => \LED_Blink_Inst.un4_r_count_5hz_cry_4\
        );

    \I__186\ : InMux
    port map (
            O => \N__2159\,
            I => \LED_Blink_Inst.un4_r_count_5hz_cry_5\
        );

    \I__185\ : InMux
    port map (
            O => \N__2156\,
            I => \LED_Blink_Inst.un4_r_count_5hz_cry_6\
        );

    \I__184\ : InMux
    port map (
            O => \N__2153\,
            I => \LED_Blink_Inst.un4_r_count_5hz_cry_7\
        );

    \IN_MUX_bfv_11_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_3_0_\
        );

    \IN_MUX_bfv_11_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \LED_Blink_Inst.un6_r_count_10hz_cry_8\,
            carryinitout => \bfn_11_4_0_\
        );

    \IN_MUX_bfv_11_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \LED_Blink_Inst.un6_r_count_10hz_cry_16\,
            carryinitout => \bfn_11_5_0_\
        );

    \IN_MUX_bfv_7_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_5_0_\
        );

    \IN_MUX_bfv_7_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \LED_Blink_Inst.un4_r_count_5hz_cry_8\,
            carryinitout => \bfn_7_6_0_\
        );

    \IN_MUX_bfv_7_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \LED_Blink_Inst.un4_r_count_5hz_cry_16\,
            carryinitout => \bfn_7_7_0_\
        );

    \IN_MUX_bfv_12_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_6_0_\
        );

    \IN_MUX_bfv_12_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \LED_Blink_Inst.un4_r_count_2hz_cry_8\,
            carryinitout => \bfn_12_7_0_\
        );

    \IN_MUX_bfv_12_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \LED_Blink_Inst.un4_r_count_2hz_cry_16\,
            carryinitout => \bfn_12_8_0_\
        );

    \IN_MUX_bfv_8_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_7_0_\
        );

    \IN_MUX_bfv_8_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \LED_Blink_Inst.un4_r_count_1hz_cry_8\,
            carryinitout => \bfn_8_8_0_\
        );

    \IN_MUX_bfv_8_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \LED_Blink_Inst.un4_r_count_1hz_cry_16\,
            carryinitout => \bfn_8_9_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \LED_Blink_Inst.un4_r_count_5hz_cry_1_c_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2391\,
            in2 => \N__2720\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_5_0_\,
            carryout => \LED_Blink_Inst.un4_r_count_5hz_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_2_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2431\,
            in2 => \_gnd_net_\,
            in3 => \N__2171\,
            lcout => \LED_Blink_Inst.r_Count_5HZZ0Z_2\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_5hz_cry_1\,
            carryout => \LED_Blink_Inst.un4_r_count_5hz_cry_2\,
            clk => \N__4428\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_3_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2296\,
            in2 => \_gnd_net_\,
            in3 => \N__2168\,
            lcout => \LED_Blink_Inst.r_Count_5HZZ0Z_3\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_5hz_cry_2\,
            carryout => \LED_Blink_Inst.un4_r_count_5hz_cry_3\,
            clk => \N__4428\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_4_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2443\,
            in2 => \_gnd_net_\,
            in3 => \N__2165\,
            lcout => \LED_Blink_Inst.r_Count_5HZZ0Z_4\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_5hz_cry_3\,
            carryout => \LED_Blink_Inst.un4_r_count_5hz_cry_4\,
            clk => \N__4428\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_RNO_0_5_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2308\,
            in2 => \_gnd_net_\,
            in3 => \N__2162\,
            lcout => \LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_5hz_cry_4\,
            carryout => \LED_Blink_Inst.un4_r_count_5hz_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_6_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2416\,
            in2 => \_gnd_net_\,
            in3 => \N__2159\,
            lcout => \LED_Blink_Inst.r_Count_5HZZ0Z_6\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_5hz_cry_5\,
            carryout => \LED_Blink_Inst.un4_r_count_5hz_cry_6\,
            clk => \N__4428\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_RNO_0_7_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2404\,
            in2 => \_gnd_net_\,
            in3 => \N__2156\,
            lcout => \LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_5hz_cry_6\,
            carryout => \LED_Blink_Inst.un4_r_count_5hz_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_RNO_0_8_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2372\,
            in2 => \_gnd_net_\,
            in3 => \N__2153\,
            lcout => \LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_5hz_cry_7\,
            carryout => \LED_Blink_Inst.un4_r_count_5hz_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_9_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2671\,
            in2 => \_gnd_net_\,
            in3 => \N__2198\,
            lcout => \LED_Blink_Inst.r_Count_5HZZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_7_6_0_\,
            carryout => \LED_Blink_Inst.un4_r_count_5hz_cry_9\,
            clk => \N__4425\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_RNO_0_10_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2464\,
            in2 => \_gnd_net_\,
            in3 => \N__2195\,
            lcout => \LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_5hz_cry_9\,
            carryout => \LED_Blink_Inst.un4_r_count_5hz_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_11_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2734\,
            in2 => \_gnd_net_\,
            in3 => \N__2192\,
            lcout => \LED_Blink_Inst.r_Count_5HZZ0Z_11\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_5hz_cry_10\,
            carryout => \LED_Blink_Inst.un4_r_count_5hz_cry_11\,
            clk => \N__4425\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_12_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2632\,
            in2 => \_gnd_net_\,
            in3 => \N__2189\,
            lcout => \LED_Blink_Inst.r_Count_5HZZ0Z_12\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_5hz_cry_11\,
            carryout => \LED_Blink_Inst.un4_r_count_5hz_cry_12\,
            clk => \N__4425\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_RNO_0_13_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2332\,
            in2 => \_gnd_net_\,
            in3 => \N__2186\,
            lcout => \LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_5hz_cry_12\,
            carryout => \LED_Blink_Inst.un4_r_count_5hz_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_14_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2659\,
            in2 => \_gnd_net_\,
            in3 => \N__2183\,
            lcout => \LED_Blink_Inst.r_Count_5HZZ0Z_14\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_5hz_cry_13\,
            carryout => \LED_Blink_Inst.un4_r_count_5hz_cry_14\,
            clk => \N__4425\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_15_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2221\,
            in2 => \_gnd_net_\,
            in3 => \N__2180\,
            lcout => \LED_Blink_Inst.r_Count_5HZZ0Z_15\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_5hz_cry_14\,
            carryout => \LED_Blink_Inst.un4_r_count_5hz_cry_15\,
            clk => \N__4425\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_16_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2644\,
            in2 => \_gnd_net_\,
            in3 => \N__2177\,
            lcout => \LED_Blink_Inst.r_Count_5HZZ0Z_16\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_5hz_cry_15\,
            carryout => \LED_Blink_Inst.un4_r_count_5hz_cry_16\,
            clk => \N__4425\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_RNO_0_17_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2683\,
            in2 => \_gnd_net_\,
            in3 => \N__2174\,
            lcout => \LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \bfn_7_7_0_\,
            carryout => \LED_Blink_Inst.un4_r_count_5hz_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_RNO_0_18_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2321\,
            in2 => \_gnd_net_\,
            in3 => \N__2276\,
            lcout => \LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_5hz_cry_17\,
            carryout => \LED_Blink_Inst.un4_r_count_5hz_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_19_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2251\,
            in2 => \_gnd_net_\,
            in3 => \N__2273\,
            lcout => \LED_Blink_Inst.r_Count_5HZZ0Z_19\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_5hz_cry_18\,
            carryout => \LED_Blink_Inst.un4_r_count_5hz_cry_19\,
            clk => \N__4423\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_20_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2242\,
            in2 => \_gnd_net_\,
            in3 => \N__2270\,
            lcout => \LED_Blink_Inst.r_Count_5HZZ0Z_20\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_5hz_cry_19\,
            carryout => \LED_Blink_Inst.un4_r_count_5hz_cry_20\,
            clk => \N__4423\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_RNO_0_21_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2233\,
            in2 => \_gnd_net_\,
            in3 => \N__2267\,
            lcout => \LED_Blink_Inst.r_Count_5HZ_RNO_0Z0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_18_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__2498\,
            in1 => \N__2264\,
            in2 => \N__2619\,
            in3 => \N__2560\,
            lcout => \LED_Blink_Inst.r_Count_5HZZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4423\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_21_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__2620\,
            in1 => \N__2499\,
            in2 => \N__2564\,
            in3 => \N__2258\,
            lcout => \LED_Blink_Inst.r_Count_5HZZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4423\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_RNIH2F11_21_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__2252\,
            in1 => \N__2243\,
            in2 => \N__2234\,
            in3 => \N__2222\,
            lcout => \LED_Blink_Inst.un1_r_count_5hz_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_7_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__2514\,
            in1 => \N__2616\,
            in2 => \N__2562\,
            in3 => \N__2210\,
            lcout => \LED_Blink_Inst.r_Count_5HZZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4433\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_5_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__2204\,
            in1 => \N__2513\,
            in2 => \N__2621\,
            in3 => \N__2555\,
            lcout => \LED_Blink_Inst.r_Count_5HZZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4433\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_RNI96LC_1_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2444\,
            in1 => \N__2432\,
            in2 => \N__2420\,
            in3 => \N__2392\,
            lcout => \LED_Blink_Inst.un1_r_count_5hz_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_RNITRA6_7_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2405\,
            in2 => \_gnd_net_\,
            in3 => \N__2371\,
            lcout => \LED_Blink_Inst.un1_r_count_5hz_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_1_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__2393\,
            in1 => \N__2719\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \LED_Blink_Inst.r_Count_5HZZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4433\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_8_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__2515\,
            in1 => \N__2617\,
            in2 => \N__2563\,
            in3 => \N__2378\,
            lcout => \LED_Blink_Inst.r_Count_5HZZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4433\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Toggle_5HZ_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__2618\,
            in1 => \N__2516\,
            in2 => \N__2356\,
            in3 => \N__2556\,
            lcout => \o_LED_2_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4433\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_0_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__2500\,
            in1 => \N__2718\,
            in2 => \N__2612\,
            in3 => \N__2548\,
            lcout => \LED_Blink_Inst.r_Count_5HZZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4429\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_13_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__2595\,
            in1 => \N__2502\,
            in2 => \N__2561\,
            in3 => \N__2339\,
            lcout => \LED_Blink_Inst.r_Count_5HZZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4429\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_RNII1D11_10_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2333\,
            in1 => \N__2465\,
            in2 => \N__2687\,
            in3 => \N__2320\,
            lcout => OPEN,
            ltout => \LED_Blink_Inst.un1_r_count_5hz_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_RNI5I2E1_3_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__2309\,
            in1 => \N__2297\,
            in2 => \N__2285\,
            in3 => \N__2282\,
            lcout => OPEN,
            ltout => \LED_Blink_Inst.un1_r_count_5hz_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_RNIE3862_11_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__2741\,
            in1 => \N__2735\,
            in2 => \N__2723\,
            in3 => \N__2717\,
            lcout => \LED_Blink_Inst.un1_r_count_5hz_19\,
            ltout => \LED_Blink_Inst.un1_r_count_5hz_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_17_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__2596\,
            in1 => \N__2503\,
            in2 => \N__2696\,
            in3 => \N__2693\,
            lcout => \LED_Blink_Inst.r_Count_5HZZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4429\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_RNI477S_9_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2672\,
            in1 => \N__2660\,
            in2 => \N__2648\,
            in3 => \N__2633\,
            lcout => \LED_Blink_Inst.un1_r_count_5hz_15\,
            ltout => \LED_Blink_Inst.un1_r_count_5hz_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_5HZ_10_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__2544\,
            in1 => \N__2501\,
            in2 => \N__2474\,
            in3 => \N__2471\,
            lcout => \LED_Blink_Inst.r_Count_5HZZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4429\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.un4_r_count_1hz_cry_1_c_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3171\,
            in2 => \N__2860\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_7_0_\,
            carryout => \LED_Blink_Inst.un4_r_count_1hz_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_2_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2821\,
            in2 => \_gnd_net_\,
            in3 => \N__2453\,
            lcout => \LED_Blink_Inst.r_Count_1HZZ0Z_2\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_1hz_cry_1\,
            carryout => \LED_Blink_Inst.un4_r_count_1hz_cry_2\,
            clk => \N__4426\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_3_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2833\,
            in2 => \_gnd_net_\,
            in3 => \N__2450\,
            lcout => \LED_Blink_Inst.r_Count_1HZZ0Z_3\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_1hz_cry_2\,
            carryout => \LED_Blink_Inst.un4_r_count_1hz_cry_3\,
            clk => \N__4426\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_4_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2872\,
            in2 => \_gnd_net_\,
            in3 => \N__2447\,
            lcout => \LED_Blink_Inst.r_Count_1HZZ0Z_4\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_1hz_cry_3\,
            carryout => \LED_Blink_Inst.un4_r_count_1hz_cry_4\,
            clk => \N__4426\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_5_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2911\,
            in2 => \_gnd_net_\,
            in3 => \N__2768\,
            lcout => \LED_Blink_Inst.r_Count_1HZZ0Z_5\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_1hz_cry_4\,
            carryout => \LED_Blink_Inst.un4_r_count_1hz_cry_5\,
            clk => \N__4426\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_6_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2899\,
            in2 => \_gnd_net_\,
            in3 => \N__2765\,
            lcout => \LED_Blink_Inst.r_Count_1HZZ0Z_6\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_1hz_cry_5\,
            carryout => \LED_Blink_Inst.un4_r_count_1hz_cry_6\,
            clk => \N__4426\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_7_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2884\,
            in2 => \_gnd_net_\,
            in3 => \N__2762\,
            lcout => \LED_Blink_Inst.r_Count_1HZZ0Z_7\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_1hz_cry_6\,
            carryout => \LED_Blink_Inst.un4_r_count_1hz_cry_7\,
            clk => \N__4426\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_RNO_0_8_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2806\,
            in2 => \_gnd_net_\,
            in3 => \N__2759\,
            lcout => \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_1hz_cry_7\,
            carryout => \LED_Blink_Inst.un4_r_count_1hz_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_RNO_0_9_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3013\,
            in2 => \_gnd_net_\,
            in3 => \N__2756\,
            lcout => \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_8_8_0_\,
            carryout => \LED_Blink_Inst.un4_r_count_1hz_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_10_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2971\,
            in2 => \_gnd_net_\,
            in3 => \N__2753\,
            lcout => \LED_Blink_Inst.r_Count_1HZZ0Z_10\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_1hz_cry_9\,
            carryout => \LED_Blink_Inst.un4_r_count_1hz_cry_10\,
            clk => \N__4422\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_RNO_0_11_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3148\,
            in2 => \_gnd_net_\,
            in3 => \N__2750\,
            lcout => \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_1hz_cry_10\,
            carryout => \LED_Blink_Inst.un4_r_count_1hz_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_RNO_0_12_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3109\,
            in2 => \_gnd_net_\,
            in3 => \N__2747\,
            lcout => \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_1hz_cry_11\,
            carryout => \LED_Blink_Inst.un4_r_count_1hz_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_13_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2986\,
            in2 => \_gnd_net_\,
            in3 => \N__2744\,
            lcout => \LED_Blink_Inst.r_Count_1HZZ0Z_13\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_1hz_cry_12\,
            carryout => \LED_Blink_Inst.un4_r_count_1hz_cry_13\,
            clk => \N__4422\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_14_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3055\,
            in2 => \_gnd_net_\,
            in3 => \N__2795\,
            lcout => \LED_Blink_Inst.r_Count_1HZZ0Z_14\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_1hz_cry_13\,
            carryout => \LED_Blink_Inst.un4_r_count_1hz_cry_14\,
            clk => \N__4422\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_15_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2956\,
            in3 => \N__2792\,
            lcout => \LED_Blink_Inst.r_Count_1HZZ0Z_15\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_1hz_cry_14\,
            carryout => \LED_Blink_Inst.un4_r_count_1hz_cry_15\,
            clk => \N__4422\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_RNO_0_16_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3031\,
            in2 => \_gnd_net_\,
            in3 => \N__2789\,
            lcout => \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_1hz_cry_15\,
            carryout => \LED_Blink_Inst.un4_r_count_1hz_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_RNO_0_17_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3199\,
            in2 => \_gnd_net_\,
            in3 => \N__2786\,
            lcout => \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \bfn_8_9_0_\,
            carryout => \LED_Blink_Inst.un4_r_count_1hz_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_RNO_0_18_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3226\,
            in2 => \_gnd_net_\,
            in3 => \N__2783\,
            lcout => \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_1hz_cry_17\,
            carryout => \LED_Blink_Inst.un4_r_count_1hz_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_19_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3085\,
            in2 => \_gnd_net_\,
            in3 => \N__2780\,
            lcout => \LED_Blink_Inst.r_Count_1HZZ0Z_19\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_1hz_cry_18\,
            carryout => \LED_Blink_Inst.un4_r_count_1hz_cry_19\,
            clk => \N__4427\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_RNO_0_20_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3239\,
            in2 => \_gnd_net_\,
            in3 => \N__2777\,
            lcout => \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_1hz_cry_19\,
            carryout => \LED_Blink_Inst.un4_r_count_1hz_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_RNO_0_21_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3214\,
            in2 => \_gnd_net_\,
            in3 => \N__2774\,
            lcout => \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_21\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_1hz_cry_20\,
            carryout => \LED_Blink_Inst.un4_r_count_1hz_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_22_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3097\,
            in2 => \_gnd_net_\,
            in3 => \N__2771\,
            lcout => \LED_Blink_Inst.r_Count_1HZZ0Z_22\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_1hz_cry_21\,
            carryout => \LED_Blink_Inst.un4_r_count_1hz_cry_22\,
            clk => \N__4427\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_RNO_0_23_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3070\,
            in2 => \_gnd_net_\,
            in3 => \N__2996\,
            lcout => OPEN,
            ltout => \LED_Blink_Inst.r_Count_1HZ_RNO_0Z0Z_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_23_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__3371\,
            in1 => \N__3283\,
            in2 => \N__2993\,
            in3 => \N__3428\,
            lcout => \LED_Blink_Inst.r_Count_1HZZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4427\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_RNI7T7T_10_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2990\,
            in1 => \N__2975\,
            in2 => \N__2960\,
            in3 => \N__2855\,
            lcout => \LED_Blink_Inst.un1_r_count_1hz_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_8_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3286\,
            in1 => \N__3422\,
            in2 => \N__3373\,
            in3 => \N__2939\,
            lcout => \LED_Blink_Inst.r_Count_1HZZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4430\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_0_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__3420\,
            in1 => \N__3284\,
            in2 => \N__3370\,
            in3 => \N__2856\,
            lcout => \LED_Blink_Inst.r_Count_1HZZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4430\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Toggle_1HZ_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__3287\,
            in1 => \N__3423\,
            in2 => \N__2929\,
            in3 => \N__3346\,
            lcout => \o_LED_4_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4430\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_RNI2VI71_4_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2912\,
            in1 => \N__2900\,
            in2 => \N__2888\,
            in3 => \N__2873\,
            lcout => \LED_Blink_Inst.un1_r_count_1hz_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_1_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__3173\,
            in1 => \_gnd_net_\,
            in2 => \N__2861\,
            in3 => \_gnd_net_\,
            lcout => \LED_Blink_Inst.r_Count_1HZZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4430\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_RNIQMI71_1_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__2834\,
            in1 => \N__2822\,
            in2 => \N__2810\,
            in3 => \N__3172\,
            lcout => \LED_Blink_Inst.un1_r_count_1hz_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_11_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__3285\,
            in1 => \N__3421\,
            in2 => \N__3158\,
            in3 => \N__3345\,
            lcout => \LED_Blink_Inst.r_Count_1HZZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4430\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_RNIH78T_11_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3110\,
            in1 => \N__3149\,
            in2 => \N__3035\,
            in3 => \N__3014\,
            lcout => OPEN,
            ltout => \LED_Blink_Inst.un1_r_count_1hz_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_RNIF0A64_11_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3188\,
            in1 => \N__3137\,
            in2 => \N__3128\,
            in3 => \N__3125\,
            lcout => \LED_Blink_Inst.un1_r_count_1hz_21\,
            ltout => \LED_Blink_Inst.un1_r_count_1hz_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_12_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3350\,
            in1 => \N__3268\,
            in2 => \N__3119\,
            in3 => \N__3116\,
            lcout => \LED_Blink_Inst.r_Count_1HZZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4424\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_RNI45SP_23_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__3098\,
            in1 => \N__3086\,
            in2 => \N__3074\,
            in3 => \N__3056\,
            lcout => \LED_Blink_Inst.un1_r_count_1hz_16\,
            ltout => \LED_Blink_Inst.un1_r_count_1hz_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_16_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3369\,
            in1 => \N__3418\,
            in2 => \N__3044\,
            in3 => \N__3041\,
            lcout => \LED_Blink_Inst.r_Count_1HZZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4424\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_9_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3419\,
            in1 => \N__3269\,
            in2 => \N__3372\,
            in3 => \N__3020\,
            lcout => \LED_Blink_Inst.r_Count_1HZZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4424\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_20_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3281\,
            in1 => \N__3426\,
            in2 => \N__3374\,
            in3 => \N__3002\,
            lcout => \LED_Blink_Inst.r_Count_1HZZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4431\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_18_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3425\,
            in1 => \N__3280\,
            in2 => \N__3377\,
            in3 => \N__3440\,
            lcout => \LED_Blink_Inst.r_Count_1HZZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4431\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_21_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3282\,
            in1 => \N__3427\,
            in2 => \N__3375\,
            in3 => \N__3434\,
            lcout => \LED_Blink_Inst.r_Count_1HZZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4431\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_17_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__3424\,
            in1 => \N__3383\,
            in2 => \N__3376\,
            in3 => \N__3279\,
            lcout => \LED_Blink_Inst.r_Count_1HZZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4431\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_1HZ_RNI23SP_17_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3238\,
            in1 => \N__3227\,
            in2 => \N__3215\,
            in3 => \N__3200\,
            lcout => \LED_Blink_Inst.un1_r_count_1hz_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.un6_r_count_10hz_cry_1_c_LC_11_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4032\,
            in2 => \N__3680\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_3_0_\,
            carryout => \LED_Blink_Inst.un6_r_count_10hz_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_2_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4045\,
            in2 => \_gnd_net_\,
            in3 => \N__3182\,
            lcout => \LED_Blink_Inst.r_Count_10HZZ0Z_2\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un6_r_count_10hz_cry_1\,
            carryout => \LED_Blink_Inst.un6_r_count_10hz_cry_2\,
            clk => \N__4443\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_3_LC_11_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3691\,
            in2 => \_gnd_net_\,
            in3 => \N__3179\,
            lcout => \LED_Blink_Inst.r_Count_10HZZ0Z_3\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un6_r_count_10hz_cry_2\,
            carryout => \LED_Blink_Inst.un6_r_count_10hz_cry_3\,
            clk => \N__4443\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_RNO_0_4_LC_11_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3658\,
            in2 => \_gnd_net_\,
            in3 => \N__3176\,
            lcout => \LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un6_r_count_10hz_cry_3\,
            carryout => \LED_Blink_Inst.un6_r_count_10hz_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_5_LC_11_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3703\,
            in2 => \_gnd_net_\,
            in3 => \N__3467\,
            lcout => \LED_Blink_Inst.r_Count_10HZZ0Z_5\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un6_r_count_10hz_cry_4\,
            carryout => \LED_Blink_Inst.un6_r_count_10hz_cry_5\,
            clk => \N__4443\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_RNO_0_6_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3641\,
            in2 => \_gnd_net_\,
            in3 => \N__3464\,
            lcout => \LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un6_r_count_10hz_cry_5\,
            carryout => \LED_Blink_Inst.un6_r_count_10hz_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_RNO_0_7_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4072\,
            in2 => \_gnd_net_\,
            in3 => \N__3461\,
            lcout => \LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un6_r_count_10hz_cry_6\,
            carryout => \LED_Blink_Inst.un6_r_count_10hz_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_8_LC_11_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4006\,
            in2 => \_gnd_net_\,
            in3 => \N__3458\,
            lcout => \LED_Blink_Inst.r_Count_10HZZ0Z_8\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un6_r_count_10hz_cry_7\,
            carryout => \LED_Blink_Inst.un6_r_count_10hz_cry_8\,
            clk => \N__4443\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_RNO_0_9_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3961\,
            in2 => \_gnd_net_\,
            in3 => \N__3455\,
            lcout => \LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_11_4_0_\,
            carryout => \LED_Blink_Inst.un6_r_count_10hz_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_10_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3994\,
            in2 => \_gnd_net_\,
            in3 => \N__3452\,
            lcout => \LED_Blink_Inst.r_Count_10HZZ0Z_10\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un6_r_count_10hz_cry_9\,
            carryout => \LED_Blink_Inst.un6_r_count_10hz_cry_10\,
            clk => \N__4441\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_11_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3577\,
            in2 => \_gnd_net_\,
            in3 => \N__3449\,
            lcout => \LED_Blink_Inst.r_Count_10HZZ0Z_11\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un6_r_count_10hz_cry_10\,
            carryout => \LED_Blink_Inst.un6_r_count_10hz_cry_11\,
            clk => \N__4441\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_RNO_0_12_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4084\,
            in2 => \_gnd_net_\,
            in3 => \N__3446\,
            lcout => \LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un6_r_count_10hz_cry_11\,
            carryout => \LED_Blink_Inst.un6_r_count_10hz_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_13_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3616\,
            in2 => \_gnd_net_\,
            in3 => \N__3443\,
            lcout => \LED_Blink_Inst.r_Count_10HZZ0Z_13\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un6_r_count_10hz_cry_12\,
            carryout => \LED_Blink_Inst.un6_r_count_10hz_cry_13\,
            clk => \N__4441\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_14_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3589\,
            in2 => \_gnd_net_\,
            in3 => \N__3521\,
            lcout => \LED_Blink_Inst.r_Count_10HZZ0Z_14\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un6_r_count_10hz_cry_13\,
            carryout => \LED_Blink_Inst.un6_r_count_10hz_cry_14\,
            clk => \N__4441\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_15_LC_11_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3604\,
            in2 => \_gnd_net_\,
            in3 => \N__3518\,
            lcout => \LED_Blink_Inst.r_Count_10HZZ0Z_15\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un6_r_count_10hz_cry_14\,
            carryout => \LED_Blink_Inst.un6_r_count_10hz_cry_15\,
            clk => \N__4441\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_RNO_0_16_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4058\,
            in2 => \_gnd_net_\,
            in3 => \N__3515\,
            lcout => \LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un6_r_count_10hz_cry_15\,
            carryout => \LED_Blink_Inst.un6_r_count_10hz_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_RNO_0_17_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3529\,
            in2 => \_gnd_net_\,
            in3 => \N__3512\,
            lcout => \LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \bfn_11_5_0_\,
            carryout => \LED_Blink_Inst.un6_r_count_10hz_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_18_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3475\,
            in2 => \_gnd_net_\,
            in3 => \N__3509\,
            lcout => \LED_Blink_Inst.r_Count_10HZZ0Z_18\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un6_r_count_10hz_cry_17\,
            carryout => \LED_Blink_Inst.un6_r_count_10hz_cry_18\,
            clk => \N__4439\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_19_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3484\,
            in2 => \_gnd_net_\,
            in3 => \N__3506\,
            lcout => \LED_Blink_Inst.r_Count_10HZZ0Z_19\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un6_r_count_10hz_cry_18\,
            carryout => \LED_Blink_Inst.un6_r_count_10hz_cry_19\,
            clk => \N__4439\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_RNO_0_20_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3497\,
            in2 => \_gnd_net_\,
            in3 => \N__3503\,
            lcout => OPEN,
            ltout => \LED_Blink_Inst.r_Count_10HZ_RNO_0Z0Z_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_20_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__3832\,
            in1 => \N__3945\,
            in2 => \N__3500\,
            in3 => \N__3879\,
            lcout => \LED_Blink_Inst.r_Count_10HZZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4439\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_RNI9JA61_20_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__3530\,
            in1 => \N__3496\,
            in2 => \N__3488\,
            in3 => \N__3476\,
            lcout => \LED_Blink_Inst.un1_r_count_10hz_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_17_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__3878\,
            in1 => \N__3536\,
            in2 => \N__3950\,
            in3 => \N__3833\,
            lcout => \LED_Blink_Inst.r_Count_10HZZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4439\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_1_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3763\,
            in2 => \_gnd_net_\,
            in3 => \N__3782\,
            lcout => \LED_Blink_Inst.r_Count_2HZZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4436\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_RNIPIKC_6_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__4175\,
            in1 => \N__4190\,
            in2 => \_gnd_net_\,
            in3 => \N__3761\,
            lcout => \LED_Blink_Inst.un1_r_count_2hz_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_RNIR7RG_1_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3725\,
            in1 => \N__3781\,
            in2 => \N__4208\,
            in3 => \N__3740\,
            lcout => \LED_Blink_Inst.un1_r_count_2hz_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_11_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__4578\,
            in1 => \N__4097\,
            in2 => \N__4528\,
            in3 => \N__4643\,
            lcout => \LED_Blink_Inst.r_Count_2HZZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4435\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_0_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__3762\,
            in1 => \N__4641\,
            in2 => \N__4529\,
            in3 => \N__4580\,
            lcout => \LED_Blink_Inst.r_Count_2HZZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4435\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_4_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__4579\,
            in1 => \N__4524\,
            in2 => \N__4220\,
            in3 => \N__4644\,
            lcout => \LED_Blink_Inst.r_Count_2HZZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4435\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_RNI009U_4_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4136\,
            in1 => \N__4157\,
            in2 => \N__4112\,
            in3 => \N__4232\,
            lcout => \LED_Blink_Inst.un1_r_count_2hz_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_9_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__4519\,
            in1 => \N__4645\,
            in2 => \N__4591\,
            in3 => \N__4145\,
            lcout => \LED_Blink_Inst.r_Count_2HZZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4435\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_10_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__4642\,
            in1 => \N__4520\,
            in2 => \N__4124\,
            in3 => \N__4584\,
            lcout => \LED_Blink_Inst.r_Count_2HZZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4435\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_16_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__4638\,
            in1 => \N__4573\,
            in2 => \N__4298\,
            in3 => \N__4513\,
            lcout => \LED_Blink_Inst.r_Count_2HZZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4432\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_20_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__4511\,
            in1 => \N__4640\,
            in2 => \N__4590\,
            in3 => \N__4241\,
            lcout => \LED_Blink_Inst.r_Count_2HZZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4432\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_19_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__4639\,
            in1 => \N__4574\,
            in2 => \N__4265\,
            in3 => \N__4514\,
            lcout => \LED_Blink_Inst.r_Count_2HZZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4432\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_RNI7QMB1_12_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4310\,
            in1 => \N__4334\,
            in2 => \N__4682\,
            in3 => \N__4367\,
            lcout => OPEN,
            ltout => \LED_Blink_Inst.un1_r_count_2hz_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_RNIRKF73_1_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3566\,
            in1 => \N__3560\,
            in2 => \N__3554\,
            in3 => \N__3551\,
            lcout => \LED_Blink_Inst.un1_r_count_2hz_20\,
            ltout => \LED_Blink_Inst.un1_r_count_2hz_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_14_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__4571\,
            in1 => \N__4637\,
            in2 => \N__3545\,
            in3 => \N__4322\,
            lcout => \LED_Blink_Inst.r_Count_2HZZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4432\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_12_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__4636\,
            in1 => \N__4572\,
            in2 => \N__4355\,
            in3 => \N__4512\,
            lcout => \LED_Blink_Inst.r_Count_2HZZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4432\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_RNI9UOB1_22_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4661\,
            in1 => \N__4253\,
            in2 => \N__4757\,
            in3 => \N__4277\,
            lcout => \LED_Blink_Inst.un1_r_count_2hz_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_0_LC_12_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__3678\,
            in1 => \N__3885\,
            in2 => \N__3948\,
            in3 => \N__3830\,
            lcout => \LED_Blink_Inst.r_Count_10HZZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4445\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_7_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3829\,
            in1 => \N__3940\,
            in2 => \N__3893\,
            in3 => \N__3542\,
            lcout => \LED_Blink_Inst.r_Count_10HZZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4445\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_4_LC_12_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__3884\,
            in1 => \N__3710\,
            in2 => \N__3949\,
            in3 => \N__3831\,
            lcout => \LED_Blink_Inst.r_Count_10HZZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4445\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_RNI1U1B_3_LC_12_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__3704\,
            in1 => \N__3692\,
            in2 => \_gnd_net_\,
            in3 => \N__3677\,
            lcout => \LED_Blink_Inst.un1_r_count_10hz_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_1_LC_12_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__3679\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4034\,
            lcout => \LED_Blink_Inst.r_Count_10HZZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4445\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_RNIG3C7_4_LC_12_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3659\,
            in2 => \_gnd_net_\,
            in3 => \N__3640\,
            lcout => \LED_Blink_Inst.un1_r_count_10hz_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_6_LC_12_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3828\,
            in1 => \N__3939\,
            in2 => \N__3892\,
            in3 => \N__3647\,
            lcout => \LED_Blink_Inst.r_Count_10HZZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4445\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_16_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__3881\,
            in1 => \N__3629\,
            in2 => \N__3947\,
            in3 => \N__3835\,
            lcout => \LED_Blink_Inst.r_Count_10HZZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4444\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_12_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__3880\,
            in1 => \N__3623\,
            in2 => \N__3946\,
            in3 => \N__3834\,
            lcout => \LED_Blink_Inst.r_Count_10HZZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4444\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_RNIT5961_11_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3617\,
            in1 => \N__3605\,
            in2 => \N__3593\,
            in3 => \N__3578\,
            lcout => \LED_Blink_Inst.un1_r_count_10hz_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_RNI6UGQ_7_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4085\,
            in1 => \N__3962\,
            in2 => \N__4073\,
            in3 => \N__4057\,
            lcout => OPEN,
            ltout => \LED_Blink_Inst.un1_r_count_10hz_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_RNIVT891_1_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__4046\,
            in1 => \N__4033\,
            in2 => \N__4016\,
            in3 => \N__4013\,
            lcout => OPEN,
            ltout => \LED_Blink_Inst.un1_r_count_10hz_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_RNIV6J12_8_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__4007\,
            in1 => \N__3995\,
            in2 => \N__3983\,
            in3 => \N__3980\,
            lcout => \LED_Blink_Inst.un1_r_count_10hz_18\,
            ltout => \LED_Blink_Inst.un1_r_count_10hz_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_10HZ_9_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__3883\,
            in1 => \N__3971\,
            in2 => \N__3965\,
            in3 => \N__3932\,
            lcout => \LED_Blink_Inst.r_Count_10HZZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4444\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Toggle_10HZ_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__3941\,
            in1 => \N__3882\,
            in2 => \N__3797\,
            in3 => \N__3836\,
            lcout => \o_LED_1_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4442\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.un4_r_count_2hz_cry_1_c_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3780\,
            in2 => \N__3764\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_6_0_\,
            carryout => \LED_Blink_Inst.un4_r_count_2hz_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_2_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3739\,
            in2 => \_gnd_net_\,
            in3 => \N__3728\,
            lcout => \LED_Blink_Inst.r_Count_2HZZ0Z_2\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_2hz_cry_1\,
            carryout => \LED_Blink_Inst.un4_r_count_2hz_cry_2\,
            clk => \N__4440\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_3_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3724\,
            in2 => \_gnd_net_\,
            in3 => \N__3713\,
            lcout => \LED_Blink_Inst.r_Count_2HZZ0Z_3\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_2hz_cry_2\,
            carryout => \LED_Blink_Inst.un4_r_count_2hz_cry_3\,
            clk => \N__4440\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_RNO_0_4_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4231\,
            in2 => \_gnd_net_\,
            in3 => \N__4211\,
            lcout => \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_2hz_cry_3\,
            carryout => \LED_Blink_Inst.un4_r_count_2hz_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_5_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4204\,
            in2 => \_gnd_net_\,
            in3 => \N__4193\,
            lcout => \LED_Blink_Inst.r_Count_2HZZ0Z_5\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_2hz_cry_4\,
            carryout => \LED_Blink_Inst.un4_r_count_2hz_cry_5\,
            clk => \N__4440\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_6_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4189\,
            in2 => \_gnd_net_\,
            in3 => \N__4178\,
            lcout => \LED_Blink_Inst.r_Count_2HZZ0Z_6\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_2hz_cry_5\,
            carryout => \LED_Blink_Inst.un4_r_count_2hz_cry_6\,
            clk => \N__4440\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_7_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4174\,
            in2 => \_gnd_net_\,
            in3 => \N__4163\,
            lcout => \LED_Blink_Inst.r_Count_2HZZ0Z_7\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_2hz_cry_6\,
            carryout => \LED_Blink_Inst.un4_r_count_2hz_cry_7\,
            clk => \N__4440\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_8_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4702\,
            in2 => \_gnd_net_\,
            in3 => \N__4160\,
            lcout => \LED_Blink_Inst.r_Count_2HZZ0Z_8\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_2hz_cry_7\,
            carryout => \LED_Blink_Inst.un4_r_count_2hz_cry_8\,
            clk => \N__4440\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_RNO_0_9_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4156\,
            in2 => \_gnd_net_\,
            in3 => \N__4139\,
            lcout => \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_12_7_0_\,
            carryout => \LED_Blink_Inst.un4_r_count_2hz_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_RNO_0_10_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4135\,
            in2 => \_gnd_net_\,
            in3 => \N__4115\,
            lcout => \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_2hz_cry_9\,
            carryout => \LED_Blink_Inst.un4_r_count_2hz_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_RNO_0_11_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4108\,
            in2 => \_gnd_net_\,
            in3 => \N__4088\,
            lcout => \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_2hz_cry_10\,
            carryout => \LED_Blink_Inst.un4_r_count_2hz_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_RNO_0_12_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4366\,
            in2 => \_gnd_net_\,
            in3 => \N__4340\,
            lcout => \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_2hz_cry_11\,
            carryout => \LED_Blink_Inst.un4_r_count_2hz_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_13_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4729\,
            in2 => \_gnd_net_\,
            in3 => \N__4337\,
            lcout => \LED_Blink_Inst.r_Count_2HZZ0Z_13\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_2hz_cry_12\,
            carryout => \LED_Blink_Inst.un4_r_count_2hz_cry_13\,
            clk => \N__4437\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_RNO_0_14_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4333\,
            in2 => \_gnd_net_\,
            in3 => \N__4316\,
            lcout => \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_2hz_cry_13\,
            carryout => \LED_Blink_Inst.un4_r_count_2hz_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_15_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4741\,
            in2 => \_gnd_net_\,
            in3 => \N__4313\,
            lcout => \LED_Blink_Inst.r_Count_2HZZ0Z_15\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_2hz_cry_14\,
            carryout => \LED_Blink_Inst.un4_r_count_2hz_cry_15\,
            clk => \N__4437\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_RNO_0_16_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4309\,
            in2 => \_gnd_net_\,
            in3 => \N__4286\,
            lcout => \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_2hz_cry_15\,
            carryout => \LED_Blink_Inst.un4_r_count_2hz_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_RNO_0_17_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4678\,
            in2 => \_gnd_net_\,
            in3 => \N__4283\,
            lcout => \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \bfn_12_8_0_\,
            carryout => \LED_Blink_Inst.un4_r_count_2hz_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_RNO_0_18_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4660\,
            in2 => \_gnd_net_\,
            in3 => \N__4280\,
            lcout => \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_2hz_cry_17\,
            carryout => \LED_Blink_Inst.un4_r_count_2hz_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_RNO_0_19_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4276\,
            in2 => \_gnd_net_\,
            in3 => \N__4256\,
            lcout => \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_2hz_cry_18\,
            carryout => \LED_Blink_Inst.un4_r_count_2hz_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_RNO_0_20_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4252\,
            in2 => \_gnd_net_\,
            in3 => \N__4235\,
            lcout => \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_2hz_cry_19\,
            carryout => \LED_Blink_Inst.un4_r_count_2hz_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_21_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4714\,
            in2 => \_gnd_net_\,
            in3 => \N__4766\,
            lcout => \LED_Blink_Inst.r_Count_2HZZ0Z_21\,
            ltout => OPEN,
            carryin => \LED_Blink_Inst.un4_r_count_2hz_cry_20\,
            carryout => \LED_Blink_Inst.un4_r_count_2hz_cry_21\,
            clk => \N__4434\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_RNO_0_22_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4756\,
            in2 => \_gnd_net_\,
            in3 => \N__4763\,
            lcout => OPEN,
            ltout => \LED_Blink_Inst.r_Count_2HZ_RNO_0Z0Z_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_22_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__4570\,
            in1 => \N__4646\,
            in2 => \N__4760\,
            in3 => \N__4518\,
            lcout => \LED_Blink_Inst.r_Count_2HZZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4434\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_RNILV051_8_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4742\,
            in1 => \N__4730\,
            in2 => \N__4718\,
            in3 => \N__4706\,
            lcout => \LED_Blink_Inst.un1_r_count_2hz_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_17_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__4647\,
            in1 => \N__4586\,
            in2 => \N__4691\,
            in3 => \N__4516\,
            lcout => \LED_Blink_Inst.r_Count_2HZZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4438\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Count_2HZ_18_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__4515\,
            in1 => \N__4648\,
            in2 => \N__4592\,
            in3 => \N__4667\,
            lcout => \LED_Blink_Inst.r_Count_2HZZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4438\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_Blink_Inst.r_Toggle_2HZ_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__4649\,
            in1 => \N__4585\,
            in2 => \N__4462\,
            in3 => \N__4517\,
            lcout => \o_LED_3_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4438\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
